CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
640 80 30 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
47
9 2-In NOR~
219 1062 361 0 1 22
0 0
0
0 0 608 90
6 74LS02
-21 -24 21 -16
4 U11B
-289 -267 -261 -259
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
7376 0 0
2
44300.9 0
0
9 2-In NOR~
219 838 365 0 1 22
0 0
0
0 0 608 90
6 74LS02
-21 -24 21 -16
4 U11A
-53 -285 -25 -277
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
9156 0 0
2
44300.9 0
0
14 Logic Display~
6 1059 128 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5776 0 0
2
44300.9 1
0
14 Logic Display~
6 1104 128 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7207 0 0
2
44300.9 0
0
13 Logic Switch~
5 1175 232 0 1 11
0 12
0
0 0 21344 90
2 0V
11 0 25 8
2 S5
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4459 0 0
2
44300.9 2
0
13 Logic Switch~
5 1214 232 0 1 11
0 10
0
0 0 21344 90
2 0V
11 0 25 8
2 S4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3760 0 0
2
44300.9 1
0
13 Logic Switch~
5 1254 235 0 1 11
0 11
0
0 0 21344 90
2 0V
11 0 25 8
2 S3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
754 0 0
2
44300.9 0
0
9 Inverter~
13 872 355 0 2 22
0 17 25
0
0 0 608 90
5 74F04
-18 -19 17 -11
3 U3E
-158 -311 -137 -303
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
9767 0 0
2
44300.9 13
0
9 Inverter~
13 1098 359 0 2 22
0 16 21
0
0 0 608 90
5 74F04
-18 -19 17 -11
3 U3D
-296 -311 -275 -303
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
7978 0 0
2
44300.9 12
0
9 2-In AND~
219 911 355 0 3 22
0 17 15 24
0
0 0 608 90
5 74F08
-18 -24 17 -16
3 U4D
-188 -308 -167 -300
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3142 0 0
2
44300.9 11
0
9 2-In AND~
219 1132 357 0 3 22
0 16 14 20
0
0 0 608 90
5 74F08
-18 -24 17 -16
3 U4C
-358 -293 -337 -285
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3284 0 0
2
44300.9 10
0
8 2-In OR~
219 943 360 0 3 22
0 17 15 23
0
0 0 608 90
5 74F32
-18 -24 17 -16
4 U10B
-261 -310 -233 -302
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
659 0 0
2
44300.9 9
0
8 2-In OR~
219 1165 360 0 3 22
0 16 14 19
0
0 0 608 90
5 74F32
-18 -24 17 -16
4 U10A
-412 -322 -384 -314
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
3800 0 0
2
44300.9 8
0
9 2-In XOR~
219 982 359 0 3 22
0 17 15 22
0
0 0 608 90
5 74F86
-18 -24 17 -16
3 U6D
-260 -311 -239 -303
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
6792 0 0
2
44300.9 7
0
9 2-In XOR~
219 1205 362 0 3 22
0 16 14 18
0
0 0 608 90
5 74F86
-18 -24 17 -16
3 U6C
-421 -314 -400 -306
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3701 0 0
2
44300.9 6
0
5 7401~
219 1018 355 0 3 22
0 17 15 9
0
0 0 608 90
6 74LS01
-21 -24 21 -16
3 U7D
-325 -291 -304 -283
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 2 3 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
6316 0 0
2
44300.9 5
0
5 7401~
219 1242 356 0 3 22
0 16 14 8
0
0 0 608 90
6 74LS01
-21 -24 21 -16
3 U7C
-495 -291 -474 -283
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 2 3 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
8734 0 0
2
44300.9 4
0
13 Logic Switch~
5 952 461 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21344 90
2 5V
-6 21 8 29
2 A3
-6 33 8 41
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7988 0 0
2
44300.9 3
0
13 Logic Switch~
5 997 464 0 1 11
0 16
0
0 0 21344 90
2 0V
-6 17 8 25
2 A2
-5 32 9 40
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3217 0 0
2
44300.9 2
0
13 Logic Switch~
5 1130 456 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21344 90
2 5V
-8 17 6 25
2 B3
-5 33 9 41
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3965 0 0
2
44300.9 1
0
13 Logic Switch~
5 1171 462 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21344 90
2 5V
-5 16 9 24
2 B2
-3 29 11 37
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8239 0 0
2
44300.9 0
0
7 74LS151
20 1095 243 0 1 29
0 0
0
0 0 4832 90
6 74F151
-21 -60 21 -52
2 U9
-313 -231 -299 -223
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 0 0 0 0
1 U
828 0 0
2
44300.9 0
0
7 74LS151
20 978 245 0 1 29
0 0
0
0 0 4832 90
6 74F151
-21 -60 21 -52
2 U8
-207 -233 -193 -225
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 0 0 0 0
1 U
6187 0 0
2
44300.9 0
0
13 Logic Switch~
5 175 100 0 1 11
0 11
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 S0
-6 -37 8 -29
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7107 0 0
2
5.89981e-315 0
0
13 Logic Switch~
5 135 97 0 1 11
0 10
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 S1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6433 0 0
2
5.89981e-315 0
0
13 Logic Switch~
5 96 97 0 1 11
0 12
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 S2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8559 0 0
2
5.89981e-315 0
0
13 Logic Switch~
5 467 416 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21344 90
2 5V
-5 16 9 24
2 B0
-3 29 11 37
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3674 0 0
2
44300.9 0
0
13 Logic Switch~
5 426 410 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21344 90
2 5V
-8 17 6 25
2 B1
-5 33 9 41
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5697 0 0
2
44300.9 1
0
13 Logic Switch~
5 293 418 0 1 11
0 16
0
0 0 21344 90
2 0V
-6 17 8 25
2 A0
-5 32 9 40
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3805 0 0
2
44300.9 2
0
13 Logic Switch~
5 248 415 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21344 90
2 5V
-6 21 8 29
2 A1
-6 33 8 41
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5219 0 0
2
44300.9 3
0
14 Logic Display~
6 380 81 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3795 0 0
2
5.89981e-315 0
0
14 Logic Display~
6 325 82 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3637 0 0
2
5.89981e-315 0
0
8 2-In OR~
219 377 141 0 3 22
0 6 4 2
0
0 0 608 90
5 74F32
-18 -24 17 -16
3 U5D
-258 -310 -237 -302
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3226 0 0
2
5.89981e-315 0
0
8 2-In OR~
219 321 138 0 3 22
0 7 5 3
0
0 0 608 90
5 74F32
-18 -24 17 -16
3 U5C
-258 -310 -237 -302
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
6966 0 0
2
5.89981e-315 0
0
9 Inverter~
13 129 255 0 2 22
0 12 13
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U3C
-148 -186 -127 -178
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
9796 0 0
2
5.89981e-315 0
0
5 7401~
219 553 309 0 3 22
0 16 14 8
0
0 0 608 90
6 74LS01
-21 -24 21 -16
3 U7B
-495 -291 -474 -283
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 2 3 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
5952 0 0
2
44300.9 4
0
5 7401~
219 316 308 0 3 22
0 17 15 9
0
0 0 608 90
6 74LS01
-21 -24 21 -16
3 U7A
-325 -291 -304 -283
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 2 3 1 2 3 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3649 0 0
2
44300.9 5
0
9 2-In XOR~
219 509 317 0 3 22
0 16 14 18
0
0 0 608 90
5 74F86
-18 -24 17 -16
3 U6B
-421 -314 -400 -306
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3716 0 0
2
44300.9 6
0
9 2-In XOR~
219 278 313 0 3 22
0 17 15 22
0
0 0 608 90
5 74F86
-18 -24 17 -16
3 U6A
-260 -311 -239 -303
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
4797 0 0
2
44300.9 7
0
8 2-In OR~
219 471 316 0 3 22
0 16 14 19
0
0 0 608 90
5 74F32
-18 -24 17 -16
3 U5B
-409 -322 -388 -314
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
4681 0 0
2
44300.9 8
0
8 2-In OR~
219 239 314 0 3 22
0 17 15 23
0
0 0 608 90
5 74F32
-18 -24 17 -16
3 U5A
-258 -310 -237 -302
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9730 0 0
2
44300.9 9
0
9 2-In AND~
219 440 312 0 3 22
0 16 14 20
0
0 0 608 90
5 74F08
-18 -24 17 -16
3 U4B
-358 -293 -337 -285
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
9874 0 0
2
44300.9 10
0
9 2-In AND~
219 207 309 0 3 22
0 17 15 24
0
0 0 608 90
5 74F08
-18 -24 17 -16
3 U4A
-188 -308 -167 -300
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
364 0 0
2
44300.9 11
0
9 Inverter~
13 405 312 0 2 22
0 16 21
0
0 0 608 90
5 74F04
-18 -19 17 -11
3 U3B
-296 -311 -275 -303
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3656 0 0
2
44300.9 12
0
9 Inverter~
13 168 309 0 2 22
0 17 25
0
0 0 608 90
5 74F04
-18 -19 17 -11
3 U3A
-158 -311 -137 -303
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3131 0 0
2
44300.9 13
0
7 74LS257
147 450 213 0 14 29
0 13 26 9 27 8 28 29 30 31
13 5 4 32 33
0
0 0 4832 90
6 74F257
-21 -60 21 -52
2 U2
-497 -206 -483 -198
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 512 1 0 0 0
1 U
6772 0 0
2
44300.9 14
0
7 74LS153
119 314 205 0 14 29
0 25 24 23 22 10 11 21 20 19
18 12 12 7 6
0
0 0 4832 90
6 74F153
-21 -60 21 -52
2 U1
-216 -212 -202 -204
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 0 1 0 0 0
1 U
9557 0 0
2
44300.9 15
0
86
2 0 0 0 0 0 0 1 0 0 30 3
1077 380
1077 425
1140 425
1 0 0 0 0 0 0 1 0 0 44 3
1059 380
1059 405
1101 405
2 0 0 0 0 16 0 2 0 0 35 4
853 384
853 430
920 430
920 431
1 0 0 0 0 0 0 2 0 0 43 4
835 384
835 400
875 400
875 401
3 3 0 0 0 0 0 1 22 0 0 4
1068 328
1068 326
1092 326
1092 275
3 3 0 0 0 0 0 2 23 0 0 4
844 332
844 297
975 297
975 277
1 13 0 0 0 0 0 4 22 0 0 4
1104 146
1104 169
1128 169
1128 211
1 13 0 0 0 0 0 3 23 0 0 4
1059 146
1059 170
1011 170
1011 213
1 0 0 0 0 0 0 5 0 0 15 3
1176 219
1176 175
1081 175
1 0 0 0 0 0 0 6 0 0 16 4
1215 219
1215 181
1092 181
1092 180
1 0 0 0 0 0 0 7 0 0 17 3
1255 222
1255 187
1100 187
9 0 0 0 0 0 0 22 0 0 14 2
1074 205
1074 195
14 0 0 0 0 0 0 23 0 0 14 2
1020 207
1020 195
9 14 0 0 0 0 0 23 22 0 0 4
957 207
957 195
1137 195
1137 205
10 10 0 0 0 0 0 23 22 0 0 4
966 213
966 175
1083 175
1083 211
11 11 0 0 0 0 0 23 22 0 0 4
975 213
975 180
1092 180
1092 211
12 12 0 0 0 0 0 23 22 0 0 4
984 213
984 187
1101 187
1101 211
2 4 0 0 0 0 0 9 22 0 0 2
1101 341
1101 275
3 5 0 0 0 0 0 11 22 0 0 4
1131 333
1131 326
1110 326
1110 275
3 6 0 0 0 0 0 13 22 0 0 4
1168 330
1168 319
1119 319
1119 275
3 7 0 0 0 0 0 15 22 0 0 4
1208 332
1208 313
1128 313
1128 275
3 8 0 0 0 0 0 17 22 0 0 4
1244 329
1244 307
1137 307
1137 275
4 2 0 0 0 0 0 23 8 0 0 4
984 277
984 304
875 304
875 337
5 3 0 0 0 0 0 23 10 0 0 4
993 277
993 312
910 312
910 331
6 3 0 0 0 0 0 23 12 0 0 4
1002 277
1002 318
946 318
946 330
7 3 0 0 0 0 0 23 14 0 0 4
1011 277
1011 325
985 325
985 329
8 3 0 0 0 0 0 23 16 0 0 2
1020 277
1020 328
2 0 14 0 0 0 0 15 0 0 31 2
1217 381
1217 424
2 0 14 0 0 0 0 13 0 0 31 4
1177 376
1177 409
1176 409
1176 424
2 0 14 0 0 0 0 11 0 0 31 3
1140 378
1140 425
1157 425
1 2 14 0 0 0 0 21 17 0 0 5
1172 449
1157 449
1157 424
1253 424
1253 380
2 0 15 0 0 0 0 16 0 0 35 4
1029 379
1029 411
1031 411
1031 431
2 0 15 0 0 0 0 14 0 0 35 4
994 378
994 411
993 411
993 431
2 0 15 0 0 0 0 12 0 0 35 2
955 376
955 431
1 2 15 0 0 0 0 20 10 0 0 4
1131 443
1131 431
919 431
919 376
1 0 16 0 0 0 0 11 0 0 39 4
1122 378
1122 392
1121 392
1121 405
1 0 16 0 0 0 0 13 0 0 39 2
1159 376
1159 405
1 0 16 0 0 0 0 15 0 0 39 2
1199 381
1199 405
0 1 16 0 0 0 0 0 17 44 0 3
1112 405
1235 405
1235 380
1 0 17 0 0 0 0 14 0 0 43 2
976 378
976 401
1 0 17 0 0 0 0 12 0 0 43 2
937 376
937 401
1 0 17 0 0 0 0 10 0 0 43 2
901 376
901 401
0 1 17 0 0 0 0 0 16 45 0 3
875 401
1011 401
1011 379
1 1 16 0 0 0 0 19 9 0 0 6
998 451
998 441
1112 441
1112 405
1101 405
1101 377
1 1 17 0 0 0 0 18 8 0 0 4
953 448
953 442
875 442
875 373
1 3 2 0 0 12416 0 31 33 0 0 4
380 99
380 96
380 96
380 111
1 3 3 0 0 12416 0 32 34 0 0 4
325 100
325 99
324 99
324 108
2 12 4 0 0 8320 0 33 46 0 0 4
389 157
389 171
445 171
445 180
2 11 5 0 0 8320 0 34 46 0 0 4
333 154
333 163
427 163
427 180
1 14 6 0 0 8320 0 33 47 0 0 4
371 157
371 167
342 167
342 178
1 13 7 0 0 8320 0 34 47 0 0 4
315 154
315 166
297 166
297 178
3 5 8 0 0 8320 0 36 46 0 0 4
555 282
555 267
445 267
445 244
3 3 9 0 0 8320 0 37 46 0 0 4
318 281
318 269
427 269
427 244
5 1 10 0 0 8320 0 47 25 0 0 4
315 242
315 244
135 244
135 109
1 6 11 0 0 8320 0 24 47 0 0 4
175 112
175 249
324 249
324 242
11 0 12 0 0 0 0 47 0 0 57 2
279 172
279 172
12 0 12 0 0 4224 0 47 0 0 60 2
360 172
96 172
1 0 13 0 0 8192 0 46 0 0 59 3
409 244
410 244
410 254
2 10 13 0 0 4224 0 35 46 0 0 5
150 255
410 255
410 254
490 254
490 250
1 1 12 0 0 0 0 26 35 0 0 3
96 109
96 255
114 255
2 0 14 0 0 4096 0 38 0 0 64 2
521 336
521 378
2 0 14 0 0 4096 0 40 0 0 64 2
483 332
483 378
2 0 14 0 0 0 0 42 0 0 64 3
448 333
448 379
453 379
1 2 14 0 0 12416 0 27 36 0 0 5
468 403
453 403
453 378
564 378
564 333
2 0 15 0 0 4096 0 37 0 0 68 2
327 332
327 380
2 0 15 0 0 0 0 39 0 0 68 4
290 332
290 365
289 365
289 380
2 0 15 0 0 4096 0 41 0 0 68 2
251 330
251 380
1 2 15 0 0 8320 0 28 43 0 0 4
427 397
427 380
215 380
215 330
1 0 16 0 0 4096 0 42 0 0 72 2
430 333
430 359
1 0 16 0 0 4096 0 40 0 0 72 2
465 332
465 359
1 0 16 0 0 0 0 38 0 0 72 2
503 336
503 359
0 1 16 0 0 4224 0 0 36 77 0 3
408 359
546 359
546 333
1 0 17 0 0 4096 0 39 0 0 76 2
272 332
272 355
1 0 17 0 0 4096 0 41 0 0 76 2
233 330
233 355
1 0 17 0 0 0 0 43 0 0 76 2
197 330
197 355
0 1 17 0 0 4224 0 0 37 78 0 3
171 355
309 355
309 332
1 1 16 0 0 0 0 29 44 0 0 4
294 405
294 395
408 395
408 330
1 1 17 0 0 0 0 30 45 0 0 4
249 402
249 396
171 396
171 327
3 10 18 0 0 8320 0 38 47 0 0 4
512 287
512 274
360 274
360 242
3 9 19 0 0 8320 0 40 47 0 0 4
474 286
474 280
351 280
351 242
3 8 20 0 0 8320 0 42 47 0 0 4
439 288
439 286
342 286
342 242
2 7 21 0 0 8320 0 44 47 0 0 4
408 294
408 289
333 289
333 242
3 4 22 0 0 12416 0 39 47 0 0 4
281 283
281 282
306 282
306 242
3 3 23 0 0 8320 0 41 47 0 0 4
242 284
242 274
297 274
297 242
3 2 24 0 0 8320 0 43 47 0 0 4
206 285
206 267
288 267
288 242
2 1 25 0 0 8320 0 45 47 0 0 4
171 291
171 261
279 261
279 242
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
556 126 741 147
564 133 732 148
21 S2  S1  S0  Operation
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
567 158 696 179
575 165 687 180
14 0  0  0   X-OR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
567 179 680 200
575 186 671 201
12 0  0  1   OR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
567 200 682 221
576 207 672 222
12 0  1  0  AND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
566 221 689 242
575 227 679 242
13 0  1  1   NOT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
568 239 697 260
576 246 688 261
14 1  0  0   NAND
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
