CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 150 30 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
33
13 Logic Switch~
5 118 226 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-31 -4 -17 4
2 V3
1092 479 1106 487
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89969e-315 5.26354e-315
0
13 Logic Switch~
5 120 200 0 1 11
0 2
0
0 0 21344 0
2 0V
-34 -3 -20 5
2 V4
1099 463 1113 471
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89969e-315 0
0
13 Logic Switch~
5 633 929 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89969e-315 0
0
13 Logic Switch~
5 70 819 0 1 11
0 10
0
0 0 21344 0
2 0V
-31 -4 -17 4
2 V6
1092 479 1106 487
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89969e-315 5.32571e-315
0
13 Logic Switch~
5 72 793 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-34 -3 -20 5
2 V5
1099 463 1113 471
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.89969e-315 5.30499e-315
0
13 Logic Switch~
5 767 393 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.89969e-315 0
0
13 Logic Switch~
5 767 271 0 1 11
0 21
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
5.89969e-315 0
0
9 2-In AND~
219 421 269 0 3 22
0 3 2 8
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
7361 0 0
2
5.89969e-315 5.40342e-315
0
8 2-In OR~
219 411 348 0 3 22
0 3 2 7
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
4747 0 0
2
5.89969e-315 5.39824e-315
0
9 2-In NOR~
219 416 516 0 3 22
0 3 2 5
0
0 0 608 0
6 74LS02
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
972 0 0
2
5.89969e-315 5.39306e-315
0
14 Logic Display~
6 560 265 0 1 2
10 8
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L3
-8 -14 6 -6
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
5.89969e-315 5.38788e-315
0
10 2-In NAND~
219 427 430 0 3 22
0 3 2 6
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9998 0 0
2
5.89969e-315 5.37752e-315
0
14 Logic Display~
6 560 344 0 1 2
10 7
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L4
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
5.89969e-315 5.36716e-315
0
14 Logic Display~
6 558 426 0 1 2
10 6
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L5
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
5.89969e-315 5.3568e-315
0
14 Logic Display~
6 562 512 0 1 2
10 5
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L6
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
5.89969e-315 5.34643e-315
0
14 Logic Display~
6 564 600 0 1 2
10 4
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L8
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
5.89969e-315 5.32571e-315
0
9 2-In XOR~
219 416 604 0 3 22
0 3 2 4
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
5616 0 0
2
5.89969e-315 5.30499e-315
0
14 Logic Display~
6 885 925 0 1 2
10 11
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L13
-8 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
5.89969e-315 5.30499e-315
0
9 Inverter~
13 743 929 0 2 22
0 12 11
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U3D
-7 -17 14 -9
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
317 0 0
2
5.89969e-315 5.26354e-315
0
9 2-In AND~
219 371 839 0 3 22
0 10 9 17
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3108 0 0
2
5.89969e-315 5.40342e-315
0
8 2-In OR~
219 363 916 0 3 22
0 10 9 16
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U2B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
4299 0 0
2
5.89969e-315 5.39824e-315
0
9 2-In NOR~
219 367 1066 0 3 22
0 10 9 14
0
0 0 608 0
6 74LS02
-21 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
9672 0 0
2
5.89969e-315 5.39306e-315
0
14 Logic Display~
6 510 835 0 1 2
10 17
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L12
-11 -14 10 -6
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
5.89969e-315 5.38788e-315
0
10 2-In NAND~
219 371 989 0 3 22
0 10 9 15
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
6369 0 0
2
5.89969e-315 5.37752e-315
0
14 Logic Display~
6 510 912 0 1 2
10 16
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L11
-8 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
5.89969e-315 5.36716e-315
0
14 Logic Display~
6 509 985 0 1 2
10 15
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L10
-8 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
5.89969e-315 5.3568e-315
0
14 Logic Display~
6 513 1062 0 1 2
10 14
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L9
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
5.89969e-315 5.34643e-315
0
14 Logic Display~
6 516 1139 0 1 2
10 13
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L7
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
5.89969e-315 5.26354e-315
0
9 2-In XOR~
219 368 1143 0 3 22
0 10 9 13
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U6B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
961 0 0
2
5.89969e-315 0
0
9 Inverter~
13 862 393 0 2 22
0 19 18
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
3178 0 0
2
5.89969e-315 5.30499e-315
0
14 Logic Display~
6 1021 389 0 1 2
10 18
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
5.89969e-315 5.26354e-315
0
9 Inverter~
13 877 272 0 2 22
0 21 20
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U3C
-7 -17 14 -9
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
3951 0 0
2
5.89969e-315 5.30499e-315
0
14 Logic Display~
6 1019 268 0 1 2
10 20
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8885 0 0
2
5.89969e-315 5.26354e-315
0
36
2 0 2 0 0 4096 0 10 0 0 9 2
403 525
150 525
1 0 3 0 0 4096 0 10 0 0 10 2
403 507
130 507
2 0 2 0 0 0 0 12 0 0 9 2
403 439
150 439
1 0 3 0 0 0 0 12 0 0 10 2
403 421
130 421
2 0 2 0 0 0 0 9 0 0 9 2
398 357
150 357
1 0 3 0 0 0 0 9 0 0 10 2
398 339
130 339
2 0 2 0 0 0 0 8 0 0 9 2
397 278
150 278
1 0 3 0 0 0 0 8 0 0 10 2
397 260
130 260
1 2 2 0 0 8320 0 2 17 0 0 4
132 200
150 200
150 613
400 613
1 1 3 0 0 4224 0 1 17 0 0 3
130 226
130 595
400 595
1 3 4 0 0 4224 0 16 17 0 0 2
548 604
449 604
1 3 5 0 0 4224 0 15 10 0 0 2
546 516
455 516
1 3 6 0 0 4224 0 14 12 0 0 2
542 430
454 430
1 3 7 0 0 4224 0 13 9 0 0 2
544 348
444 348
1 3 8 0 0 4224 0 11 8 0 0 2
544 269
442 269
2 0 9 0 0 4096 0 22 0 0 25 2
354 1075
101 1075
1 0 10 0 0 4096 0 22 0 0 24 2
354 1057
82 1057
2 0 9 0 0 0 0 24 0 0 25 2
347 998
101 998
1 0 10 0 0 0 0 24 0 0 24 2
347 980
82 980
2 0 9 0 0 0 0 21 0 0 25 2
350 925
101 925
1 0 10 0 0 0 0 21 0 0 24 2
350 907
82 907
2 0 9 0 0 0 0 20 0 0 25 2
347 848
101 848
1 0 10 0 0 0 0 20 0 0 24 2
347 830
82 830
1 1 10 0 0 4224 0 4 29 0 0 3
82 819
82 1134
352 1134
1 2 9 0 0 8320 0 5 29 0 0 4
84 793
101 793
101 1152
352 1152
2 1 11 0 0 4224 0 19 18 0 0 2
764 929
869 929
1 1 12 0 0 4224 0 3 19 0 0 2
645 929
728 929
1 3 13 0 0 4224 0 28 29 0 0 2
500 1143
401 1143
1 3 14 0 0 4224 0 27 22 0 0 2
497 1066
406 1066
1 3 15 0 0 4224 0 26 24 0 0 2
493 989
398 989
1 3 16 0 0 4224 0 25 21 0 0 2
494 916
396 916
1 3 17 0 0 4224 0 23 20 0 0 2
494 839
392 839
1 2 18 0 0 4224 0 31 30 0 0 2
1005 393
883 393
1 1 19 0 0 4224 0 6 30 0 0 2
779 393
847 393
1 2 20 0 0 4224 0 33 32 0 0 2
1003 272
898 272
1 1 21 0 0 8320 0 7 32 0 0 3
779 271
779 272
862 272
85
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
266 198 323 219
274 205 314 220
5 B = 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
266 176 323 197
274 183 314 198
5 A = 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
214 175 275 199
224 183 264 199
5 Input
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
275 352 340 373
283 359 331 374
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
384 366 459 387
393 373 449 388
7 OR Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
718 141 817 163
727 148 807 164
10 INPUT  A B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
722 169 807 193
732 177 796 193
8 OUTPUT X
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
924 245 991 267
933 253 981 269
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
791 246 858 268
800 254 848 270
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
747 276 856 300
757 284 845 300
11 INPUT A = 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
824 458 909 482
834 466 898 482
8 NOT Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
888 275 995 297
897 282 985 298
11 Output X =1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
910 359 977 381
919 367 967 383
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
781 355 848 377
790 363 838 379
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
754 399 863 423
764 407 852 423
11 INPUT A = 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
897 399 1004 421
906 406 994 422
11 Output X =0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
331 1164 416 1188
341 1172 405 1188
8 XOR Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
220 1112 287 1134
229 1120 277 1136
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
217 1144 284 1166
226 1152 274 1168
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
421 1114 488 1136
430 1122 478 1138
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
420 1038 487 1060
429 1045 477 1061
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
223 1068 290 1090
232 1075 280 1091
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
417 962 484 984
426 970 474 986
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
214 957 281 979
223 964 271 980
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
415 887 482 909
424 894 472 910
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
216 882 283 904
225 890 273 906
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
403 814 470 836
412 821 460 837
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
217 804 284 826
226 811 274 827
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
220 1034 287 1056
229 1042 277 1058
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
213 990 280 1012
222 998 270 1014
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
213 917 280 939
222 925 270 941
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
214 841 281 863
223 849 271 865
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
325 852 410 876
335 859 399 875
8 AND Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
329 1077 414 1101
339 1085 403 1101
8 NOR Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
325 1002 418 1026
335 1010 407 1026
9 NAND Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
330 928 407 952
340 936 396 952
7 OR Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
657 904 724 926
666 912 714 928
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
790 903 857 925
799 911 847 927
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
119 805 146 826
128 812 136 827
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
123 846 150 867
132 853 140 868
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
115 885 140 906
123 892 131 907
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
123 925 150 946
132 932 140 947
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
116 955 141 976
124 962 132 977
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
117 993 142 1014
125 999 133 1014
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
115 1033 140 1054
123 1040 131 1055
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
115 1075 140 1096
123 1082 131 1097
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
119 1115 146 1136
128 1122 136 1137
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
121 1150 146 1171
129 1157 137 1172
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
643 933 670 954
652 939 660 954
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
468 574 535 595
477 581 525 596
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
273 570 338 591
281 576 329 591
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
58 186 91 207
66 192 82 207
2 B=
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
58 210 93 231
67 217 83 232
2 A=
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
211 614 236 635
219 621 227 636
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
213 516 238 537
221 523 229 538
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
214 433 239 454
222 440 230 455
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
212 351 237 372
220 358 228 373
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
211 569 238 590
220 575 228 590
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
213 486 240 507
222 492 230 507
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
212 399 239 420
221 405 229 420
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
210 317 237 338
219 323 227 338
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
212 272 237 293
220 279 228 294
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
209 237 236 258
218 243 226 258
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
381 614 466 638
391 622 455 638
8 XOR Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
268 614 335 636
277 622 325 638
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
465 488 532 510
474 495 522 511
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
274 519 341 541
283 526 331 542
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
463 400 530 422
472 408 520 424
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
280 395 347 417
289 402 337 418
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
463 322 530 344
472 329 520 345
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
275 310 342 332
284 318 332 334
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
457 244 524 266
466 251 514 267
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
275 236 342 258
284 243 332 259
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
277 482 344 504
286 490 334 506
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
280 434 347 456
289 442 337 458
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
274 273 341 295
283 281 331 297
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
381 282 466 306
391 289 455 305
8 AND Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
383 530 468 554
393 538 457 554
8 NOR Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
378 446 471 470
388 454 460 470
9 NAND Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
605 210 674 232
615 217 663 233
6 Output
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
613 257 670 278
621 263 661 278
5 X = 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
617 418 674 439
625 425 665 440
5 X = 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
608 333 667 354
617 340 657 355
5 X = 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
621 500 678 521
629 507 669 522
5 X = 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
615 586 674 607
624 593 664 608
5 X = 1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
