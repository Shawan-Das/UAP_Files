CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
950 580 1 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.326954 0.500000
176 502 1364 707
42991634 0
0
6 Title:
5 Name:
0
0
0
51
13 Logic Switch~
5 1171 991 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3932 0 0
2
44283.6 0
0
13 Logic Switch~
5 1166 949 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5288 0 0
2
44283.6 0
0
13 Logic Switch~
5 1251 763 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4934 0 0
2
44283.6 0
0
13 Logic Switch~
5 1255 617 0 1 11
0 59
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 1 0 -1 0
1 V
5987 0 0
2
44283.6 0
0
13 Logic Switch~
5 1179 481 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7737 0 0
2
44283.6 0
0
13 Logic Switch~
5 1286 307 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4200 0 0
2
5.89978e-315 0
0
5 SCOPE
12 1453 670 0 1 11
0 2
0
0 0 57584 0
3 TP3
-11 -4 10 4
3 U19
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
5780 0 0
2
44283.7 0
0
5 SCOPE
12 1408 670 0 1 11
0 3
0
0 0 57584 0
3 TP2
-11 -4 10 4
3 U18
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
6490 0 0
2
44283.7 0
0
5 SCOPE
12 1370 670 0 1 11
0 4
0
0 0 57584 0
3 TP1
-11 -4 10 4
3 U17
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
8663 0 0
2
44283.7 0
0
14 Logic Display~
6 1396 934 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
318 0 0
2
44283.6 0
0
5 4027~
219 1340 995 0 7 32
0 60 6 8 5 61 62 7
0
0 0 4720 0
4 4027
7 -60 35 -52
4 U16A
-32 -61 -4 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 7 0
1 U
348 0 0
2
44283.6 0
0
5 4027~
219 1343 842 0 7 32
0 63 2 8 2 64 65 4
0
0 0 4720 0
4 4027
7 -60 35 -52
4 U15B
-32 -61 -4 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 6 0
1 U
8551 0 0
2
44283.6 7
0
5 4027~
219 1447 840 0 7 32
0 10 9 8 9 66 67 3
0
0 0 4720 0
4 4027
7 -60 35 -52
4 U15A
13 -59 41 -51
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 6 0
1 U
7295 0 0
2
44283.6 6
0
5 4027~
219 1570 840 0 7 32
0 68 3 8 3 69 70 2
0
0 0 4720 0
4 4027
7 -60 35 -52
4 U14B
12 -62 40 -54
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 5 0
1 U
9900 0 0
2
44283.6 5
0
7 Pulser~
4 1190 807 0 10 12
0 8 71 8 72 0 0 5 5 1
8
0
0 0 4656 0
0
2 V8
-4 -27 10 -19
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8725 0 0
2
44283.6 4
0
14 Logic Display~
6 1617 703 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
366 0 0
2
44283.6 3
0
14 Logic Display~
6 1642 702 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5762 0 0
2
44283.6 2
0
14 Logic Display~
6 1668 702 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4943 0 0
2
44283.6 1
0
14 Logic Display~
6 1596 420 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3435 0 0
2
44283.6 2
0
14 Logic Display~
6 1570 420 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8705 0 0
2
44283.6 1
0
14 Logic Display~
6 1545 421 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4331 0 0
2
44283.6 0
0
7 Pulser~
4 1118 525 0 10 12
0 16 73 16 74 0 0 5 5 1
8
0
0 0 4656 0
0
2 V4
-4 -27 10 -19
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
787 0 0
2
44283.6 0
0
5 4027~
219 1498 558 0 7 32
0 75 12 16 12 76 77 13
0
0 0 4720 0
4 4027
7 -60 35 -52
4 U14A
12 -62 40 -54
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 5 0
1 U
3655 0 0
2
44283.6 0
0
5 4027~
219 1375 558 0 7 32
0 15 14 16 14 78 79 12
0
0 0 4720 0
4 4027
7 -60 35 -52
4 U13B
13 -59 41 -51
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 4 0
1 U
6682 0 0
2
44283.6 0
0
5 4027~
219 1271 560 0 7 32
0 80 14 16 14 81 82 11
0
0 0 4720 0
4 4027
7 -60 35 -52
4 U13A
-32 -61 -4 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 4 0
1 U
582 0 0
2
44283.6 0
0
12 Hex Display~
7 1516 168 0 18 19
10 18 17 83 84 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
6 DISP10
-21 -38 21 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
3125 0 0
2
5.89978e-315 0
0
5 4027~
219 1508 341 0 7 32
0 22 20 17 20 21 85 18
0
0 0 4720 0
4 4027
7 -60 35 -52
4 U12B
23 -61 51 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 3 0
1 U
5466 0 0
2
5.89978e-315 0
0
5 4027~
219 1387 342 0 7 32
0 22 20 19 20 21 86 17
0
0 0 4720 0
4 4027
7 -60 35 -52
4 U12A
23 -61 51 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 3 0
1 U
52 0 0
2
5.89978e-315 0
0
7 Pulser~
4 1091 212 0 10 12
0 19 87 19 88 0 0 5 5 1
8
0
0 0 4656 0
0
2 V1
-4 -27 10 -19
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3898 0 0
2
44283.6 0
0
12 Hex Display~
7 1299 123 0 18 19
10 25 24 23 89 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP9
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
9413 0 0
2
44283.6 1
0
7 74LS293
154 1259 202 0 8 17
0 23 23 90 19 23 24 25 91
0
0 0 4848 0
7 74LS293
-24 -35 25 -27
3 U11
-11 -36 10 -28
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 512 1 0 0 0
1 U
8576 0 0
2
44283.6 2
0
12 Hex Display~
7 562 68 0 18 19
10 33 32 34 31 0 0 0 0 0
0 1 1 1 0 0 0 0 7
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP8
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
622 0 0
2
44283.6 3
0
7 74LS293
154 680 240 0 8 17
0 31 32 26 33 31 34 32 33
0
0 0 4848 90
7 74LS293
-24 -35 25 -27
3 U10
-440 -188 -419 -180
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 0 1 0 0 0
1 U
9152 0 0
2
44283.6 4
0
7 74LS293
154 627 240 0 8 17
0 27 28 31 30 27 29 28 30
0
0 0 4848 90
7 74LS293
-24 -35 25 -27
2 U9
-627 -226 -613 -218
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 0 1 0 0 0
1 U
783 0 0
2
44283.6 5
0
12 Hex Display~
7 531 68 0 18 19
10 30 28 29 27 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP7
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4262 0 0
2
44283.6 6
0
12 Hex Display~
7 463 70 0 16 19
10 39 38 40 36 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP6
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6121 0 0
2
44283.6 7
0
7 74LS293
154 541 239 0 8 17
0 36 38 27 39 36 40 38 39
0
0 0 4848 90
7 74LS293
-24 -35 25 -27
2 U8
-541 -220 -527 -212
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 0 1 0 0 0
1 U
3879 0 0
2
44283.6 8
0
7 74LS293
154 488 239 0 8 17
0 35 37 92 36 35 37 41 93
0
0 0 4848 90
7 74LS293
-24 -35 25 -27
2 U7
-485 -220 -471 -212
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 512 1 0 0 0
1 U
7345 0 0
2
44283.6 9
0
12 Hex Display~
7 432 70 0 16 19
10 41 37 35 94 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP5
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
3198 0 0
2
44283.6 10
0
12 Hex Display~
7 255 74 0 16 19
10 55 52 54 51 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9849 0 0
2
44283.6 11
0
7 74LS293
154 246 240 0 8 17
0 49 49 44 55 51 54 52 55
0
0 0 4848 90
7 74LS293
-24 -35 25 -27
2 U6
-924 -218 -910 -210
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 0 1 0 0 0
1 U
479 0 0
2
44283.6 12
0
7 74LS293
154 194 240 0 8 17
0 50 50 95 51 57 53 58 96
0
0 0 4848 90
7 74LS293
-24 -35 25 -27
2 U5
-885 -218 -871 -210
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 512 1 0 0 0
1 U
3905 0 0
2
44283.6 13
0
12 Hex Display~
7 224 74 0 16 19
10 58 53 57 97 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP4
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
4394 0 0
2
44283.6 14
0
9 2-In AND~
219 140 286 0 3 22
0 53 54 50
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
4391 0 0
2
44283.6 15
0
8 2-In OR~
219 223 319 0 3 22
0 50 56 49
0
0 0 624 90
5 74F32
-18 -24 17 -16
3 U4A
-123 -2 -102 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3681 0 0
2
44283.6 16
0
9 2-In AND~
219 269 340 0 3 22
0 51 52 56
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U3A
-14 -38 7 -30
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
6466 0 0
2
44283.6 17
0
12 Hex Display~
7 325 73 0 16 19
10 48 43 44 98 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
5230 0 0
2
44283.6 18
0
7 74LS293
154 347 240 0 8 17
0 44 43 99 42 44 43 48 100
0
0 0 4848 90
7 74LS293
-24 -35 25 -27
2 U1
-349 -214 -335 -206
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 512 1 0 0 0
1 U
8324 0 0
2
44283.6 19
0
7 74LS293
154 400 240 0 8 17
0 42 45 35 46 42 47 45 46
0
0 0 4848 90
7 74LS293
-24 -35 25 -27
2 U2
-437 -188 -423 -180
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 0 1 0 0 0
1 U
3445 0 0
2
44283.6 20
0
12 Hex Display~
7 358 73 0 16 19
10 46 45 47 42 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
7543 0 0
2
44283.6 21
0
7 Pulser~
4 484 321 0 10 12
0 101 102 26 103 0 0 5 5 1
8
0
0 0 4656 0
0
2 V2
-4 -27 10 -19
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6187 0 0
2
44283.6 22
0
116
0 1 2 0 0 4096 0 0 7 9 0 2
1453 738
1453 682
0 1 3 0 0 4096 0 0 8 11 0 4
1481 804
1481 690
1408 690
1408 682
0 1 4 0 0 4096 0 0 9 13 0 4
1378 806
1378 690
1370 690
1370 682
0 4 2 0 0 0 0 0 12 9 0 3
1311 806
1311 824
1319 824
1 4 5 0 0 4224 0 1 11 0 0 4
1183 991
1308 991
1308 977
1316 977
1 2 6 0 0 4224 0 2 11 0 0 4
1178 949
1308 949
1308 959
1316 959
7 1 7 0 0 4224 0 11 10 0 0 3
1364 959
1396 959
1396 952
0 3 8 0 0 4096 0 0 11 18 0 3
1236 815
1236 968
1316 968
0 2 2 0 0 4224 0 0 12 12 0 4
1617 738
1311 738
1311 806
1319 806
1 0 3 0 0 8320 0 17 0 0 11 4
1642 720
1642 778
1495 778
1495 804
7 0 3 0 0 0 0 13 0 0 20 2
1471 804
1538 804
7 1 2 0 0 128 0 14 16 0 0 3
1594 804
1617 804
1617 721
7 1 4 0 0 12416 0 12 18 0 0 5
1367 806
1409 806
1409 753
1668 753
1668 720
1 0 9 0 0 4224 0 3 0 0 21 4
1263 763
1400 763
1400 814
1415 814
1 0 10 0 0 4224 0 13 0 0 0 2
1447 783
1447 777
3 0 8 0 0 0 0 13 0 0 17 3
1423 813
1419 813
1419 859
0 3 8 0 0 8320 0 0 14 18 0 5
1255 815
1255 859
1533 859
1533 813
1546 813
3 0 8 0 0 0 0 12 0 0 19 2
1319 815
1225 815
1 3 8 0 0 0 0 15 15 0 0 6
1166 798
1153 798
1153 830
1225 830
1225 798
1214 798
2 4 3 0 0 0 0 14 14 0 0 4
1546 804
1538 804
1538 822
1546 822
2 4 9 0 0 0 0 13 13 0 0 4
1423 804
1415 804
1415 822
1423 822
7 1 11 0 0 12416 0 25 19 0 0 5
1295 524
1313 524
1313 488
1596 488
1596 438
0 1 12 0 0 8320 0 0 20 32 0 4
1431 522
1431 475
1570 475
1570 438
7 1 13 0 0 8320 0 23 21 0 0 3
1522 522
1545 522
1545 439
1 0 14 0 0 4096 0 5 0 0 31 2
1191 481
1230 481
1 0 15 0 0 4224 0 24 0 0 0 2
1375 501
1375 495
3 0 16 0 0 8192 0 24 0 0 28 3
1351 531
1347 531
1347 577
0 3 16 0 0 8320 0 0 23 29 0 5
1183 533
1183 577
1461 577
1461 531
1474 531
3 0 16 0 0 0 0 25 0 0 30 2
1247 533
1153 533
1 3 16 0 0 0 0 22 22 0 0 6
1094 516
1081 516
1081 548
1153 548
1153 516
1142 516
0 0 14 0 0 12416 0 0 0 35 34 6
1343 532
1333 532
1333 466
1230 466
1230 524
1239 524
7 0 12 0 0 0 0 24 0 0 33 2
1399 522
1466 522
2 4 12 0 0 0 0 23 23 0 0 4
1474 522
1466 522
1466 540
1474 540
2 4 14 0 0 0 0 25 25 0 0 4
1247 524
1239 524
1239 542
1247 542
2 4 14 0 0 0 0 24 24 0 0 4
1351 522
1343 522
1343 540
1351 540
0 2 17 0 0 4224 0 0 26 43 0 4
1441 305
1441 200
1519 200
1519 192
7 1 18 0 0 8320 0 27 26 0 0 5
1532 305
1542 305
1542 200
1525 200
1525 192
0 3 19 0 0 8320 0 0 28 48 0 5
1162 220
1162 318
1355 318
1355 315
1363 315
1 0 20 0 0 4096 0 6 0 0 42 2
1298 307
1346 307
0 0 20 0 0 8320 0 0 0 42 41 5
1346 324
1346 349
1458 349
1458 323
1463 323
2 4 20 0 0 0 0 27 27 0 0 4
1484 305
1463 305
1463 323
1484 323
2 4 20 0 0 0 0 28 28 0 0 4
1363 306
1346 306
1346 324
1363 324
7 3 17 0 0 0 0 28 27 0 0 5
1411 306
1411 305
1442 305
1442 314
1484 314
5 5 21 0 0 8320 0 28 27 0 0 4
1387 348
1387 355
1508 355
1508 347
1 1 22 0 0 8320 0 28 27 0 0 4
1387 285
1387 276
1508 276
1508 284
0 2 23 0 0 8192 0 0 31 47 0 3
1206 192
1206 202
1227 202
0 1 23 0 0 8320 0 0 31 50 0 5
1291 193
1291 158
1206 158
1206 193
1227 193
4 0 19 0 0 0 0 31 0 0 49 2
1221 220
1126 220
1 3 19 0 0 0 0 29 29 0 0 6
1067 203
1054 203
1054 235
1126 235
1126 203
1115 203
5 3 23 0 0 0 0 31 30 0 0 3
1291 193
1296 193
1296 147
6 2 24 0 0 8320 0 31 30 0 0 3
1291 202
1302 202
1302 147
7 1 25 0 0 8320 0 31 30 0 0 3
1291 211
1308 211
1308 147
3 3 26 0 0 4224 0 51 33 0 0 3
508 312
685 312
685 276
0 3 27 0 0 4096 0 0 37 56 0 3
585 282
546 282
546 275
0 2 28 0 0 8192 0 0 34 59 0 5
632 193
592 193
592 289
623 289
623 270
5 1 27 0 0 12288 0 34 34 0 0 6
614 206
614 202
585 202
585 284
614 284
614 270
4 5 27 0 0 8320 0 35 34 0 0 4
522 92
522 129
614 129
614 206
3 6 29 0 0 8320 0 35 34 0 0 4
528 92
528 124
623 124
623 206
2 7 28 0 0 8320 0 35 34 0 0 4
534 92
534 119
632 119
632 206
1 8 30 0 0 8192 0 35 34 0 0 4
540 92
540 113
641 113
641 206
8 4 30 0 0 8320 0 34 34 0 0 6
641 206
641 202
744 202
744 289
641 289
641 276
3 0 31 0 0 8192 0 34 0 0 63 3
632 276
632 282
667 282
0 1 31 0 0 8320 0 0 33 69 0 5
667 180
717 180
717 298
667 298
667 270
0 2 32 0 0 8192 0 0 33 67 0 5
685 188
711 188
711 286
676 286
676 270
4 8 33 0 0 12288 0 33 33 0 0 6
694 276
694 280
706 280
706 198
694 198
694 206
1 8 33 0 0 8320 0 32 33 0 0 4
571 92
571 94
694 94
694 206
2 7 32 0 0 8320 0 32 33 0 0 4
565 92
565 99
685 99
685 206
3 6 34 0 0 8320 0 32 33 0 0 4
559 92
559 105
676 105
676 206
4 5 31 0 0 0 0 32 33 0 0 4
553 92
553 109
667 109
667 206
3 0 35 0 0 8192 0 49 0 0 71 3
405 276
405 280
453 280
5 1 35 0 0 12416 0 38 38 0 0 6
475 205
475 196
453 196
453 283
475 283
475 269
4 0 36 0 0 8192 0 38 0 0 74 3
502 275
502 283
528 283
6 2 37 0 0 12416 0 38 38 0 0 6
484 205
484 201
445 201
445 288
484 288
484 269
0 1 36 0 0 8320 0 0 37 80 0 5
508 179
578 179
578 297
528 297
528 269
0 2 38 0 0 8320 0 0 37 78 0 5
519 187
572 187
572 285
537 285
537 269
4 8 39 0 0 12416 0 37 37 0 0 6
555 275
555 279
567 279
567 197
555 197
555 205
1 8 39 0 0 0 0 36 37 0 0 6
472 94
472 133
523 133
523 175
555 175
555 205
2 7 38 0 0 0 0 36 37 0 0 6
466 94
466 138
519 138
519 192
546 192
546 205
3 6 40 0 0 8320 0 36 37 0 0 6
460 94
460 143
513 143
513 196
537 196
537 205
4 5 36 0 0 0 0 36 37 0 0 5
454 94
454 149
508 149
508 205
528 205
1 7 41 0 0 4224 0 39 38 0 0 4
441 94
441 156
493 156
493 205
2 6 37 0 0 0 0 39 38 0 0 4
435 94
435 162
484 162
484 205
3 5 35 0 0 0 0 39 38 0 0 4
429 94
429 170
475 170
475 205
4 0 42 0 0 8192 0 48 0 0 87 3
361 276
361 284
387 284
6 2 43 0 0 12416 0 48 48 0 0 6
343 206
343 202
304 202
304 289
343 289
343 270
0 1 44 0 0 4096 0 0 48 97 0 3
310 275
334 275
334 270
0 1 42 0 0 8320 0 0 49 93 0 5
387 180
437 180
437 298
387 298
387 270
0 2 45 0 0 8320 0 0 49 91 0 5
405 188
431 188
431 286
396 286
396 270
4 8 46 0 0 12288 0 49 49 0 0 6
414 276
414 280
426 280
426 198
414 198
414 206
1 8 46 0 0 12416 0 50 49 0 0 4
367 97
367 115
414 115
414 206
2 7 45 0 0 0 0 50 49 0 0 4
361 97
361 128
405 128
405 206
3 6 47 0 0 12416 0 50 49 0 0 4
355 97
355 139
396 139
396 206
4 5 42 0 0 0 0 50 49 0 0 4
349 97
349 150
387 150
387 206
1 7 48 0 0 4224 0 47 48 0 0 4
334 97
334 162
352 162
352 206
2 6 43 0 0 0 0 47 48 0 0 4
328 97
328 170
343 170
343 206
3 5 44 0 0 4224 0 47 48 0 0 4
322 97
322 179
334 179
334 206
5 3 44 0 0 0 0 48 41 0 0 4
334 206
310 206
310 276
251 276
1 2 49 0 0 4096 0 41 41 0 0 2
233 270
242 270
1 2 50 0 0 4096 0 42 42 0 0 2
181 270
190 270
0 1 51 0 0 8192 0 0 46 101 0 4
280 269
296 269
296 349
287 349
0 4 51 0 0 8320 0 0 42 106 0 5
233 202
280 202
280 289
208 289
208 276
0 2 52 0 0 8320 0 0 46 108 0 3
251 189
287 189
287 331
0 1 53 0 0 8320 0 0 44 115 0 4
190 183
113 183
113 277
116 277
0 2 54 0 0 4224 0 0 44 107 0 4
242 163
104 163
104 295
116 295
0 4 55 0 0 8192 0 0 41 109 0 5
260 202
275 202
275 284
260 284
260 276
4 5 51 0 0 0 0 40 41 0 0 4
246 98
246 134
233 134
233 206
3 6 54 0 0 0 0 40 41 0 0 4
252 98
252 149
242 149
242 206
2 7 52 0 0 0 0 40 41 0 0 4
258 98
258 158
251 158
251 206
1 8 55 0 0 8320 0 40 41 0 0 5
264 98
263 98
263 185
260 185
260 206
0 1 50 0 0 12288 0 0 42 113 0 4
180 286
180 287
181 287
181 270
3 1 49 0 0 4224 0 45 41 0 0 4
226 289
226 277
233 277
233 270
3 2 56 0 0 4224 0 46 45 0 0 3
242 340
235 340
235 335
3 1 50 0 0 8320 0 44 45 0 0 5
161 286
180 286
180 339
217 339
217 335
5 3 57 0 0 4224 0 42 43 0 0 4
181 206
181 117
221 117
221 98
6 2 53 0 0 0 0 42 43 0 0 4
190 206
190 123
227 123
227 98
7 1 58 0 0 4224 0 42 43 0 0 4
199 206
199 130
233 130
233 98
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
