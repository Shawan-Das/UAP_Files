CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
420 160 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
86
13 Logic Switch~
5 312 660 0 1 11
0 46
0
0 0 21360 270
2 0V
-6 -22 8 -14
2 B0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89976e-315 0
0
13 Logic Switch~
5 283 661 0 10 11
0 37 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -22 8 -14
2 B1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89976e-315 0
0
13 Logic Switch~
5 254 662 0 1 11
0 27
0
0 0 21360 270
2 0V
-6 -22 8 -14
2 B2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89976e-315 0
0
13 Logic Switch~
5 229 664 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -22 8 -14
2 B3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89976e-315 0
0
13 Logic Switch~
5 403 651 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 S0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
5.89976e-315 0
0
13 Logic Switch~
5 370 653 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 S1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
5.89976e-315 0
0
13 Logic Switch~
5 186 669 0 1 11
0 43
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.89976e-315 0
0
13 Logic Switch~
5 157 670 0 1 11
0 34
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
5.89976e-315 0
0
13 Logic Switch~
5 126 669 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4747 0 0
2
5.89976e-315 0
0
13 Logic Switch~
5 99 669 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
972 0 0
2
5.89976e-315 0
0
13 Logic Switch~
5 444 657 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-7 -20 7 -12
4 Cin1
-13 -31 15 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3472 0 0
2
5.89976e-315 0
0
13 Logic Switch~
5 548 296 0 10 11
0 55 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-34 -2 -20 6
3 Cin
-58 -3 -37 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9998 0 0
2
44264.9 0
0
13 Logic Switch~
5 546 329 0 1 11
0 53
0
0 0 21360 0
2 0V
-35 -4 -21 4
2 A0
-53 -6 -39 2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3536 0 0
2
44264.9 1
0
13 Logic Switch~
5 544 402 0 10 11
0 59 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-35 -4 -21 4
2 S0
-53 -6 -39 2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4597 0 0
2
44264.9 2
0
13 Logic Switch~
5 543 435 0 10 11
0 57 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-35 -5 -21 3
2 S1
-54 -5 -40 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3835 0 0
2
44264.9 3
0
13 Logic Switch~
5 546 368 0 10 11
0 58 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-34 -2 -20 6
2 B0
-54 -3 -40 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3670 0 0
2
44264.9 4
0
13 Logic Switch~
5 77 374 0 10 11
0 65 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-34 -2 -20 6
2 B0
-54 -3 -40 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5616 0 0
2
44264.9 5
0
13 Logic Switch~
5 74 441 0 10 11
0 64 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-35 -5 -21 3
2 S1
-54 -5 -40 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9323 0 0
2
44264.9 6
0
13 Logic Switch~
5 75 408 0 10 11
0 66 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-35 -4 -21 4
2 S0
-53 -6 -39 2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
317 0 0
2
44264.9 7
0
13 Logic Switch~
5 73 82 0 1 11
0 70
0
0 0 21360 0
2 0V
-35 -4 -21 4
1 B
-50 -6 -43 2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3108 0 0
2
44264.9 8
0
13 Logic Switch~
5 72 115 0 10 11
0 71 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-35 -5 -21 3
1 A
-51 -5 -44 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4299 0 0
2
44264.9 9
0
13 Logic Switch~
5 75 48 0 1 11
0 72
0
0 0 21360 0
2 0V
-34 -2 -20 6
3 Cin
-58 -3 -37 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9672 0 0
2
44264.9 10
0
14 Logic Display~
6 1051 662 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
5.89976e-315 0
0
14 Logic Display~
6 1088 661 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
5.89976e-315 5.39306e-315
0
9 2-In XOR~
219 794 1133 0 3 22
0 14 15 13
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U12D
1074 -372 1102 -364
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 12 0
1 U
9172 0 0
2
5.89976e-315 5.38788e-315
0
9 2-In XOR~
219 929 1106 0 3 22
0 8 13 11
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U12C
929 -333 957 -325
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
7100 0 0
2
5.89976e-315 5.37752e-315
0
9 2-In AND~
219 808 1186 0 3 22
0 15 14 16
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U13D
1058 -431 1086 -423
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 13 0
1 U
3820 0 0
2
5.89976e-315 5.36716e-315
0
9 2-In AND~
219 906 1161 0 3 22
0 13 8 12
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U13C
960 -385 988 -377
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
7678 0 0
2
5.89976e-315 5.3568e-315
0
8 2-In OR~
219 988 1170 0 3 22
0 12 16 4
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U10D
869 -400 897 -392
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
961 0 0
2
5.89976e-315 5.34643e-315
0
9 2-In AND~
219 596 1127 0 3 22
0 17 2 20
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U13B
1269 -358 1297 -350
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
3178 0 0
2
5.89976e-315 5.32571e-315
0
9 2-In AND~
219 600 1182 0 3 22
0 18 3 19
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U13A
1270 -432 1298 -424
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
3409 0 0
2
5.89976e-315 5.30499e-315
0
8 2-In OR~
219 690 1159 0 3 22
0 20 19 15
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U10C
1174 -393 1202 -385
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
3951 0 0
2
5.89976e-315 5.26354e-315
0
9 Inverter~
13 517 1156 0 2 22
0 17 18
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4F
1355 -408 1376 -400
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 4 0
1 U
8885 0 0
2
5.89976e-315 0
0
14 Logic Display~
6 1123 660 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
5.89976e-315 5.39306e-315
0
9 2-In XOR~
219 797 986 0 3 22
0 24 25 23
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U12B
1074 -372 1102 -364
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
9265 0 0
2
5.89976e-315 5.38788e-315
0
9 2-In XOR~
219 933 958 0 3 22
0 9 23 21
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U12A
929 -333 957 -325
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
9442 0 0
2
5.89976e-315 5.37752e-315
0
9 2-In AND~
219 812 1051 0 3 22
0 25 24 26
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U11D
1058 -431 1086 -423
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
9424 0 0
2
5.89976e-315 5.36716e-315
0
9 2-In AND~
219 910 1013 0 3 22
0 23 9 22
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U11C
960 -385 988 -377
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
9968 0 0
2
5.89976e-315 5.3568e-315
0
8 2-In OR~
219 992 1022 0 3 22
0 22 26 8
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U10B
869 -400 897 -392
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
9281 0 0
2
5.89976e-315 5.34643e-315
0
9 2-In AND~
219 602 989 0 3 22
0 27 2 30
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U11B
1269 -358 1297 -350
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
8464 0 0
2
5.89976e-315 5.32571e-315
0
9 2-In AND~
219 601 1049 0 3 22
0 28 3 29
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U11A
1270 -432 1298 -424
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
7168 0 0
2
5.89976e-315 5.30499e-315
0
8 2-In OR~
219 696 1020 0 3 22
0 30 29 25
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U10A
1174 -393 1202 -385
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
3171 0 0
2
5.89976e-315 5.26354e-315
0
9 Inverter~
13 519 1031 0 2 22
0 27 28
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4E
1355 -408 1376 -400
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 4 0
1 U
4139 0 0
2
5.89976e-315 0
0
14 Logic Display~
6 1150 662 0 1 2
10 31
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6435 0 0
2
5.89976e-315 5.39306e-315
0
9 2-In XOR~
219 789 840 0 3 22
0 34 35 33
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6D
1077 -372 1098 -364
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
5283 0 0
2
5.89976e-315 5.38788e-315
0
9 2-In XOR~
219 924 817 0 3 22
0 10 33 31
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6C
932 -333 953 -325
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
6874 0 0
2
5.89976e-315 5.37752e-315
0
9 2-In AND~
219 804 905 0 3 22
0 35 34 36
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U9D
1061 -431 1082 -423
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
5305 0 0
2
5.89976e-315 5.36716e-315
0
9 2-In AND~
219 902 867 0 3 22
0 33 10 32
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U9C
963 -385 984 -377
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
34 0 0
2
5.89976e-315 5.3568e-315
0
8 2-In OR~
219 984 876 0 3 22
0 32 36 9
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U8D
872 -400 893 -392
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
969 0 0
2
5.89976e-315 5.34643e-315
0
9 2-In AND~
219 594 843 0 3 22
0 37 2 40
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U9B
1272 -358 1293 -350
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
8402 0 0
2
5.89976e-315 5.32571e-315
0
9 2-In AND~
219 593 903 0 3 22
0 38 3 39
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U9A
1273 -432 1294 -424
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
3751 0 0
2
5.89976e-315 5.30499e-315
0
8 2-In OR~
219 688 874 0 3 22
0 40 39 35
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U8C
1177 -393 1198 -385
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
4292 0 0
2
5.89976e-315 5.26354e-315
0
9 Inverter~
13 511 885 0 2 22
0 37 38
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4D
1355 -408 1376 -400
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 4 0
1 U
6118 0 0
2
5.89976e-315 0
0
9 Inverter~
13 507 750 0 2 22
0 46 47
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4C
1355 -408 1376 -400
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
34 0 0
2
5.89976e-315 5.41896e-315
0
8 2-In OR~
219 684 741 0 3 22
0 49 48 44
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U8B
1177 -393 1198 -385
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
6357 0 0
2
5.89976e-315 5.41378e-315
0
9 2-In AND~
219 596 773 0 3 22
0 47 3 48
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7D
1273 -432 1294 -424
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
319 0 0
2
5.89976e-315 5.4086e-315
0
9 2-In AND~
219 596 720 0 3 22
0 46 2 49
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7C
1272 -358 1293 -350
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
3976 0 0
2
5.89976e-315 5.40342e-315
0
8 2-In OR~
219 989 751 0 3 22
0 42 45 10
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U8A
872 -400 893 -392
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
7634 0 0
2
5.89976e-315 5.39824e-315
0
9 2-In AND~
219 903 732 0 3 22
0 5 6 42
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7B
963 -385 984 -377
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
523 0 0
2
5.89976e-315 5.39306e-315
0
9 2-In AND~
219 806 778 0 3 22
0 44 43 45
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7A
1061 -431 1082 -423
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
6748 0 0
2
5.89976e-315 5.38788e-315
0
9 2-In XOR~
219 935 683 0 3 22
0 6 5 41
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6B
932 -333 953 -325
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
6901 0 0
2
5.89976e-315 5.37752e-315
0
9 2-In XOR~
219 787 696 0 3 22
0 43 44 5
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6A
1077 -372 1098 -364
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
842 0 0
2
5.89976e-315 5.36716e-315
0
14 Logic Display~
6 1180 662 0 1 2
10 41
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3277 0 0
2
5.89976e-315 5.3568e-315
0
14 Logic Display~
6 1172 338 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4212 0 0
2
44264.9 11
0
14 Logic Display~
6 1233 302 0 1 2
10 50
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4720 0 0
2
44264.9 12
0
9 2-In XOR~
219 893 383 0 3 22
0 53 54 52
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1D
1077 -372 1098 -364
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
5551 0 0
2
44264.9 13
0
9 2-In XOR~
219 1029 355 0 3 22
0 55 52 50
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1C
932 -333 953 -325
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
6986 0 0
2
44264.9 14
0
9 2-In AND~
219 908 448 0 3 22
0 54 53 56
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5D
1061 -431 1082 -423
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
8745 0 0
2
44264.9 15
0
9 2-In AND~
219 1006 410 0 3 22
0 52 55 51
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5C
963 -385 984 -377
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
9592 0 0
2
44264.9 16
0
8 2-In OR~
219 1088 419 0 3 22
0 51 56 7
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3D
872 -400 893 -392
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
8748 0 0
2
44264.9 17
0
9 2-In AND~
219 698 386 0 3 22
0 58 59 62
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5B
1272 -358 1293 -350
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
7168 0 0
2
44264.9 18
0
9 2-In AND~
219 697 446 0 3 22
0 60 57 61
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5A
1273 -432 1294 -424
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
631 0 0
2
44264.9 19
0
8 2-In OR~
219 792 417 0 3 22
0 62 61 54
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3C
1177 -393 1198 -385
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
9466 0 0
2
44264.9 20
0
9 Inverter~
13 615 428 0 2 22
0 58 60
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4B
1355 -408 1376 -400
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
3266 0 0
2
44264.9 21
0
14 Logic Display~
6 388 392 0 1 2
10 63
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7693 0 0
2
44264.9 22
0
9 Inverter~
13 146 434 0 2 22
0 65 67
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
3723 0 0
2
44264.9 23
0
8 2-In OR~
219 323 423 0 3 22
0 69 68 63
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3440 0 0
2
44264.9 24
0
9 2-In AND~
219 228 452 0 3 22
0 67 64 68
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2D
-13 -27 8 -19
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
6263 0 0
2
44264.9 25
0
9 2-In AND~
219 229 392 0 3 22
0 65 66 69
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2C
-13 -27 8 -19
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
4900 0 0
2
44264.9 26
0
8 2-In OR~
219 542 175 0 3 22
0 76 77 75
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8783 0 0
2
44264.9 27
0
14 Logic Display~
6 677 171 0 1 2
10 75
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L9
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3221 0 0
2
44264.9 28
0
14 Logic Display~
6 677 77 0 1 2
10 74
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L8
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3215 0 0
2
44264.9 29
0
9 2-In AND~
219 407 166 0 3 22
0 73 72 76
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7903 0 0
2
44264.9 30
0
9 2-In AND~
219 248 210 0 3 22
0 71 70 77
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2A
-13 -27 8 -19
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7121 0 0
2
44264.9 31
0
9 2-In XOR~
219 416 82 0 3 22
0 72 73 74
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
4484 0 0
2
44264.9 32
0
9 2-In XOR~
219 224 91 0 3 22
0 70 71 73
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
5996 0 0
2
44264.9 33
0
112
1 0 2 0 0 4096 0 5 0 0 12 2
403 663
403 729
1 0 3 0 0 4096 0 6 0 0 14 2
370 665
370 782
3 1 4 0 0 8320 0 29 23 0 0 3
1021 1170
1051 1170
1051 680
1 0 5 0 0 4096 0 59 0 0 6 3
879 723
843 723
843 696
2 0 6 0 0 8192 0 59 0 0 7 5
879 741
832 741
832 673
825 673
825 674
3 2 5 0 0 4224 0 62 61 0 0 4
820 696
907 696
907 692
919 692
1 1 6 0 0 12416 0 61 11 0 0 5
919 674
825 674
825 673
444 673
444 669
2 0 3 0 0 4096 0 51 0 0 14 2
569 912
369 912
2 0 3 0 0 4096 0 41 0 0 14 2
577 1058
369 1058
2 0 2 0 0 4096 0 40 0 0 12 2
578 998
401 998
2 0 2 0 0 0 0 50 0 0 12 2
570 852
401 852
2 2 2 0 0 8320 0 57 30 0 0 4
572 729
401 729
401 1136
572 1136
3 1 7 0 0 8320 0 70 64 0 0 3
1121 419
1172 419
1172 356
2 2 3 0 0 8320 0 56 31 0 0 4
572 782
369 782
369 1191
576 1191
1 0 8 0 0 4096 0 26 0 0 25 2
913 1097
841 1097
1 0 9 0 0 4096 0 36 0 0 40 2
917 949
845 949
1 0 10 0 0 4096 0 46 0 0 55 2
908 808
832 808
1 3 11 0 0 4224 0 24 26 0 0 3
1088 679
1088 1106
962 1106
3 1 12 0 0 4224 0 28 29 0 0 2
927 1161
975 1161
0 1 13 0 0 8192 0 0 28 27 0 3
849 1134
849 1152
882 1152
0 2 14 0 0 4096 0 0 27 22 0 3
736 1125
736 1195
784 1195
1 1 14 0 0 8320 0 10 25 0 0 7
99 681
99 1080
665 1080
665 1125
736 1125
736 1124
778 1124
0 1 15 0 0 12416 0 0 27 24 0 4
753 1159
752 1159
752 1177
784 1177
3 2 15 0 0 0 0 32 25 0 0 6
723 1159
753 1159
753 1168
753 1168
753 1142
778 1142
2 3 8 0 0 12416 0 28 39 0 0 6
882 1170
841 1170
841 1063
1029 1063
1029 1022
1025 1022
3 2 16 0 0 8320 0 27 29 0 0 5
829 1186
829 1187
932 1187
932 1179
975 1179
3 2 13 0 0 20608 0 25 26 0 0 7
827 1133
849 1133
849 1134
872 1134
872 1116
913 1116
913 1115
0 1 17 0 0 4096 0 0 33 32 0 3
476 1107
476 1156
502 1156
2 1 18 0 0 4224 0 33 31 0 0 4
538 1156
560 1156
560 1173
576 1173
3 2 19 0 0 4224 0 31 32 0 0 4
621 1182
651 1182
651 1168
677 1168
3 1 20 0 0 4224 0 30 32 0 0 4
617 1127
650 1127
650 1150
677 1150
1 1 17 0 0 4224 0 4 30 0 0 5
229 676
229 1107
564 1107
564 1118
572 1118
1 3 21 0 0 4224 0 34 36 0 0 3
1123 678
1123 958
966 958
3 1 22 0 0 4224 0 38 39 0 0 2
931 1013
979 1013
0 1 23 0 0 8192 0 0 38 42 0 3
853 986
853 1004
886 1004
0 2 24 0 0 4096 0 0 37 37 0 3
740 977
740 1060
788 1060
1 1 24 0 0 8320 0 9 35 0 0 5
126 681
126 946
669 946
669 977
781 977
0 1 25 0 0 12416 0 0 37 39 0 4
757 1020
756 1020
756 1042
788 1042
3 2 25 0 0 0 0 42 35 0 0 4
729 1020
757 1020
757 995
781 995
2 3 9 0 0 12416 0 38 49 0 0 6
886 1022
845 1022
845 915
1021 915
1021 876
1017 876
3 2 26 0 0 4224 0 37 39 0 0 4
833 1051
931 1051
931 1031
979 1031
3 2 23 0 0 4224 0 35 36 0 0 5
830 986
876 986
876 968
917 968
917 967
0 1 27 0 0 4096 0 0 43 47 0 3
480 971
480 1031
504 1031
2 1 28 0 0 4224 0 43 41 0 0 4
540 1031
564 1031
564 1040
577 1040
3 2 29 0 0 4224 0 41 42 0 0 4
622 1049
655 1049
655 1029
683 1029
3 1 30 0 0 4224 0 40 42 0 0 4
623 989
654 989
654 1011
683 1011
1 1 27 0 0 8320 0 3 40 0 0 5
254 674
254 971
568 971
568 980
578 980
1 3 31 0 0 8320 0 44 46 0 0 3
1150 680
1150 817
957 817
3 1 32 0 0 4224 0 48 49 0 0 2
923 867
971 867
0 1 33 0 0 8192 0 0 48 57 0 3
845 840
845 858
878 858
0 2 34 0 0 4096 0 0 47 52 0 3
732 831
732 914
780 914
1 1 34 0 0 8320 0 8 45 0 0 5
157 682
157 805
661 805
661 831
773 831
0 1 35 0 0 12416 0 0 47 54 0 4
749 874
748 874
748 896
780 896
3 2 35 0 0 0 0 52 45 0 0 4
721 874
749 874
749 849
773 849
2 3 10 0 0 12416 0 48 58 0 0 6
878 876
832 876
832 786
1021 786
1021 751
1022 751
3 2 36 0 0 4224 0 47 49 0 0 4
825 905
923 905
923 885
971 885
3 2 33 0 0 4224 0 45 46 0 0 5
822 840
880 840
880 825
908 825
908 826
0 1 37 0 0 4096 0 0 53 62 0 3
472 825
472 885
496 885
2 1 38 0 0 4224 0 53 51 0 0 4
532 885
556 885
556 894
569 894
3 2 39 0 0 4224 0 51 52 0 0 4
614 903
647 903
647 883
675 883
3 1 40 0 0 4224 0 50 52 0 0 4
615 843
646 843
646 865
675 865
1 1 37 0 0 8320 0 2 50 0 0 5
283 673
283 825
560 825
560 834
570 834
1 3 41 0 0 8320 0 63 61 0 0 3
1180 680
1180 683
968 683
3 1 42 0 0 12416 0 59 58 0 0 4
924 732
938 732
938 742
976 742
0 2 43 0 0 4096 0 0 60 66 0 3
724 687
724 787
782 787
1 1 43 0 0 8320 0 7 62 0 0 3
186 681
186 687
771 687
0 1 44 0 0 12288 0 0 60 68 0 4
749 741
748 741
748 769
782 769
3 2 44 0 0 8320 0 55 62 0 0 4
717 741
749 741
749 705
771 705
3 2 45 0 0 8320 0 60 58 0 0 5
827 778
827 771
922 771
922 760
976 760
0 1 46 0 0 4096 0 0 54 74 0 3
472 709
472 750
492 750
2 1 47 0 0 4224 0 54 56 0 0 4
528 750
556 750
556 764
572 764
3 2 48 0 0 4224 0 56 55 0 0 4
617 773
647 773
647 750
671 750
3 1 49 0 0 4224 0 57 55 0 0 4
617 720
646 720
646 732
671 732
1 1 46 0 0 8320 0 1 57 0 0 5
312 672
312 709
560 709
560 711
572 711
1 3 50 0 0 8320 0 65 67 0 0 3
1233 320
1233 355
1062 355
3 1 51 0 0 4224 0 69 70 0 0 2
1027 410
1075 410
0 1 52 0 0 8192 0 0 69 85 0 3
949 383
949 401
982 401
0 2 53 0 0 4096 0 0 68 79 0 3
836 374
836 457
884 457
1 1 53 0 0 4224 0 13 66 0 0 4
558 329
765 329
765 374
877 374
0 1 54 0 0 12416 0 0 68 81 0 4
853 417
852 417
852 439
884 439
3 2 54 0 0 0 0 73 66 0 0 4
825 417
853 417
853 392
877 392
2 0 55 0 0 8192 0 69 0 0 84 3
982 419
941 419
941 346
3 2 56 0 0 4240 0 68 70 0 0 4
929 448
1021 448
1021 428
1075 428
1 1 55 0 0 12416 0 12 67 0 0 4
560 296
784 296
784 346
1013 346
3 2 52 0 0 4224 0 66 67 0 0 5
926 383
972 383
972 365
1013 365
1013 364
1 2 57 0 0 12416 0 15 72 0 0 4
555 435
570 435
570 455
673 455
0 1 58 0 0 4096 0 0 74 92 0 3
576 368
576 428
600 428
1 2 59 0 0 4224 0 14 71 0 0 4
556 402
662 402
662 395
674 395
2 1 60 0 0 4224 0 74 72 0 0 4
636 428
660 428
660 437
673 437
3 2 61 0 0 4224 0 72 73 0 0 4
718 446
751 446
751 426
779 426
3 1 62 0 0 4224 0 71 73 0 0 4
719 386
750 386
750 408
779 408
1 1 58 0 0 4224 0 16 71 0 0 4
558 368
664 368
664 377
674 377
3 1 63 0 0 4224 0 77 75 0 0 3
356 423
388 423
388 410
1 2 64 0 0 12416 0 18 78 0 0 4
86 441
101 441
101 461
204 461
0 1 65 0 0 4096 0 0 76 100 0 3
107 374
107 434
131 434
1 2 66 0 0 4224 0 19 79 0 0 4
87 408
193 408
193 401
205 401
2 1 67 0 0 4224 0 76 78 0 0 4
167 434
191 434
191 443
204 443
3 2 68 0 0 4224 0 78 77 0 0 4
249 452
282 452
282 432
310 432
3 1 69 0 0 4224 0 79 77 0 0 4
250 392
281 392
281 414
310 414
1 1 65 0 0 4224 0 17 79 0 0 4
89 374
195 374
195 383
205 383
2 0 70 0 0 8320 0 84 0 0 103 3
224 219
130 219
130 82
1 0 71 0 0 8320 0 84 0 0 104 3
224 201
151 201
151 115
1 1 70 0 0 0 0 20 86 0 0 2
85 82
208 82
1 2 71 0 0 0 0 21 86 0 0 4
84 115
167 115
167 100
208 100
2 0 72 0 0 8192 0 83 0 0 111 3
383 175
309 175
309 73
1 0 73 0 0 8192 0 83 0 0 112 3
383 157
329 157
329 91
1 3 74 0 0 4224 0 82 85 0 0 4
661 81
464 81
464 82
449 82
1 3 75 0 0 4224 0 81 80 0 0 2
661 175
575 175
3 1 76 0 0 4224 0 83 80 0 0 2
428 166
529 166
3 2 77 0 0 4224 0 84 80 0 0 4
269 210
417 210
417 184
529 184
1 1 72 0 0 4224 0 22 85 0 0 4
87 48
254 48
254 73
400 73
3 2 73 0 0 4224 0 86 85 0 0 2
257 91
400 91
171
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1167 365 1228 389
1177 373 1217 389
5 Carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1189 318 1234 342
1199 326 1223 342
3 Sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
953 414 990 438
963 422 979 438
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
952 377 989 401
962 385 978 401
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1015 386 1052 410
1025 394 1041 410
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
855 452 892 476
865 460 881 476
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
857 414 886 438
867 422 875 438
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
924 421 953 445
934 429 942 445
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1119 391 1148 415
1129 399 1137 415
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1051 426 1080 450
1061 434 1069 450
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1052 385 1081 409
1062 393 1070 409
1 4
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
1060 329 1086 350
1069 337 1076 352
1 3
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
979 360 1005 381
988 368 995 383
1 2
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
978 321 1004 342
987 329 994 344
1 1
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
638 342 664 363
647 350 654 365
1 1
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
638 375 664 396
647 383 654 398
1 2
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
713 360 739 381
722 368 729 383
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
657 412 686 436
667 420 675 436
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
655 451 684 475
665 459 673 475
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
710 421 739 445
720 429 728 445
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
574 422 603 446
584 430 592 446
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
629 403 658 427
639 411 647 427
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
754 380 783 404
764 388 772 404
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
753 424 782 448
763 432 771 448
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
816 387 845 411
826 395 834 411
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
353 396 382 420
363 404 371 420
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
284 430 313 454
294 438 302 454
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
285 386 314 410
295 394 303 410
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
160 409 189 433
170 417 178 433
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
105 428 134 452
115 436 123 452
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
241 427 270 451
251 435 259 451
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
186 457 215 481
196 465 204 481
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
188 418 217 442
198 426 206 442
1 4
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
244 366 270 387
253 374 260 389
1 3
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
169 381 195 402
178 389 185 404
1 2
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
169 348 195 369
178 356 185 371
1 1
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 17
545 200 664 219
553 206 655 219
17 AB + Cin(A XOR B)
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 12
416 128 503 147
423 135 495 148
12 Cin(A XOR B)
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 15
525 56 630 75
532 63 622 76
15 A XOR B XOR Cin
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
281 184 316 203
289 191 307 204
3 A.B
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
153 215 176 235
161 221 167 235
1 B
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
156 179 177 199
163 186 169 200
1 A
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
94 60 117 80
102 66 108 80
1 B
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
94 92 115 112
101 99 107 113
1 A
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 7
251 70 308 89
258 77 300 90
7 A XOR B
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
262 50 297 70
270 57 288 71
3 Cin
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
157 58 211 81
166 65 201 80
5 Pin-1
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
177 177 231 200
186 184 221 199
5 Pin-1
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
477 144 531 167
486 151 521 166
5 Pin-1
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
163 96 217 119
172 103 207 118
5 Pin-2
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
250 87 302 110
258 94 293 109
5 Pin-3
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
351 50 403 73
359 57 394 72
5 Pin-4
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
354 86 406 109
362 93 397 108
5 Pin-5
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
442 81 494 104
450 88 485 103
5 Pin-6
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
478 179 532 202
487 186 522 201
5 Pin-2
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
573 171 625 194
581 178 616 193
5 Pin-3
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
177 214 231 237
186 221 221 236
5 Pin-2
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
275 210 327 233
283 217 318 232
5 Pin-3
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
329 135 381 158
337 142 372 157
5 Pin-4
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
328 170 380 193
336 177 371 192
5 Pin-5
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
421 160 473 183
429 167 464 182
5 Pin-6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
350 220 447 241
358 227 438 242
10 Full Adder
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
702 712 731 736
712 720 720 736
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
651 748 680 772
661 756 669 772
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
652 704 681 728
662 712 670 728
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
524 745 553 769
534 753 542 769
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
473 747 502 771
483 755 491 771
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
608 742 637 766
618 750 626 766
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
555 774 584 798
565 782 573 798
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
554 741 583 765
564 749 572 765
1 4
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
611 690 637 711
620 698 627 713
1 3
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
533 724 559 745
542 732 549 747
1 2
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
533 685 559 706
542 693 549 708
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
948 714 977 738
958 722 966 738
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
948 753 977 777
958 761 966 777
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1016 748 1045 772
1026 756 1034 772
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
823 745 852 769
833 753 841 769
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
755 741 784 765
765 749 773 765
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
752 783 789 807
762 791 778 807
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
914 706 951 730
924 714 940 730
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
853 699 890 723
863 707 879 723
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
850 734 887 758
860 742 876 758
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
848 872 885 896
858 880 874 896
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
844 833 881 857
854 841 870 857
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
911 843 948 867
921 851 937 867
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
751 909 788 933
761 917 777 933
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
753 871 782 895
763 879 771 895
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
820 878 849 902
830 886 838 902
1 8
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
534 799 560 820
543 807 550 822
1 1
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
531 827 557 848
540 835 547 850
1 2
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
609 817 635 838
618 825 625 840
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
553 869 582 893
563 877 571 893
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
551 908 580 932
561 916 569 932
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
606 878 635 902
616 886 624 902
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
857 1019 894 1043
867 1027 883 1043
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
856 980 893 1004
866 988 882 1004
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
919 989 956 1013
929 997 945 1013
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
759 1055 796 1079
769 1063 785 1079
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
761 1017 790 1041
771 1025 779 1041
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
828 1024 857 1048
838 1032 846 1048
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1022 1026 1051 1050
1032 1034 1040 1050
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
955 1029 984 1053
965 1037 973 1053
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
956 988 985 1012
966 996 974 1012
1 4
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
542 945 568 966
551 953 558 968
1 1
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
542 974 568 995
551 982 558 997
1 2
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
617 963 643 984
626 971 633 986
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
561 1015 590 1039
571 1023 579 1039
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
559 1054 588 1078
569 1062 577 1078
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
614 1024 643 1048
624 1032 632 1048
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
658 983 687 1007
668 991 676 1007
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
657 1027 686 1051
667 1035 675 1051
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
720 990 749 1014
730 998 738 1014
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
853 1165 890 1189
863 1173 879 1189
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
852 1126 889 1150
862 1134 878 1150
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
915 1137 952 1161
925 1145 941 1161
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
755 1191 792 1215
765 1199 781 1215
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
753 1153 782 1177
763 1161 771 1177
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
824 1182 853 1206
834 1190 842 1206
1 8
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
536 1078 562 1099
545 1086 552 1101
1 1
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
536 1109 562 1130
545 1117 552 1132
1 2
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
614 1101 640 1122
623 1109 630 1124
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
558 1149 587 1173
568 1157 576 1173
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
560 1188 589 1212
570 1196 578 1212
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
611 1156 640 1180
621 1164 629 1180
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1161 610 1198 634
1171 618 1187 634
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1135 611 1172 635
1145 619 1161 635
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1105 612 1142 636
1115 620 1131 636
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1069 613 1106 637
1079 621 1095 637
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
990 654 1051 678
1000 662 1040 678
5 Carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
470 879 495 903
478 887 486 903
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
523 879 548 903
531 887 539 903
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
478 1025 503 1049
486 1033 494 1049
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
532 1029 557 1053
540 1037 548 1053
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
479 1154 504 1178
487 1162 495 1178
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
529 1150 554 1174
537 1158 545 1174
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
712 845 737 869
720 853 728 869
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
649 881 674 905
657 889 665 905
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
645 839 682 863
655 847 671 863
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1015 878 1052 902
1025 886 1041 902
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
943 843 980 867
953 851 969 867
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
942 880 979 904
952 888 968 904
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
710 1131 735 1155
718 1139 726 1155
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
653 1161 678 1185
661 1169 669 1185
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
650 1124 687 1148
660 1132 676 1148
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1011 1143 1048 1167
1021 1151 1037 1167
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
942 1137 979 1161
952 1145 968 1161
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
944 1176 981 1200
954 1184 970 1200
2 13
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
750 663 776 684
759 671 766 686
1 1
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
751 703 777 724
760 711 767 726
1 2
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
811 674 837 695
820 682 827 697
1 3
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
882 647 906 668
890 655 897 670
1 4
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
885 673 909 694
893 681 900 696
1 5
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
965 657 989 678
973 665 980 680
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
811 814 836 838
819 822 827 838
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
743 806 780 830
753 814 769 830
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
754 844 779 868
762 852 770 868
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
956 792 993 816
966 800 982 816
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
868 784 905 808
878 792 894 808
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
879 818 916 842
889 826 905 842
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
755 947 784 971
765 955 773 971
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
759 990 788 1014
769 998 777 1014
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
818 954 847 978
828 962 836 978
1 3
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
882 924 906 945
890 932 897 947
1 4
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
883 963 907 984
891 971 898 986
1 5
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
964 932 988 953
972 940 979 955
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
753 1099 782 1123
763 1107 771 1123
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
754 1133 783 1157
764 1141 772 1157
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
816 1104 845 1128
826 1112 834 1128
1 3
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
878 1072 902 1093
886 1080 893 1095
1 4
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
879 1111 903 1132
887 1119 894 1134
1 5
-12 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
960 1080 984 1101
968 1088 975 1103
1 6
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
