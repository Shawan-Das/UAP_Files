CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 90 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
33
13 Logic Switch~
5 72 512 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89968e-315 0
0
13 Logic Switch~
5 69 585 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89968e-315 0
0
14 Logic Display~
6 1085 267 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3124 0 0
2
5.89968e-315 0
0
14 Logic Display~
6 1084 182 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3421 0 0
2
5.89968e-315 0
0
14 Logic Display~
6 876 81 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.89968e-315 0
0
14 Logic Display~
6 1038 550 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
5.89968e-315 0
0
14 Logic Display~
6 946 617 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
5.89968e-315 0
0
10 2-In XNOR~
219 481 691 0 3 22
0 13 12 6
0
0 0 624 0
4 4077
-7 -24 21 -16
3 U5D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 5 0
1 U
7361 0 0
2
5.89968e-315 0
0
10 2-In XNOR~
219 646 114 0 3 22
0 9 2 8
0
0 0 624 0
4 4077
-7 -24 21 -16
3 U5C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
4747 0 0
2
5.89968e-315 0
0
10 2-In XNOR~
219 449 303 0 3 22
0 11 12 3
0
0 0 624 0
4 4077
-7 -24 21 -16
3 U5B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
972 0 0
2
5.89968e-315 0
0
9 2-In AND~
219 766 571 0 3 22
0 7 6 10
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U9D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
3472 0 0
2
5.89968e-315 0
0
9 2-In AND~
219 1011 198 0 3 22
0 15 16 4
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
9998 0 0
2
5.89968e-315 0
0
9 2-In AND~
219 272 207 0 3 22
0 2 13 11
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
3536 0 0
2
5.89968e-315 0
0
9 2-In AND~
219 199 111 0 3 22
0 13 2 18
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
4597 0 0
2
5.89968e-315 0
0
9 2-In XOR~
219 773 475 0 3 22
0 3 14 22
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U8C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 8 0
1 U
3835 0 0
2
5.89968e-315 0
0
9 2-In XOR~
219 747 205 0 3 22
0 15 17 16
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U8B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
3670 0 0
2
5.89968e-315 0
0
9 2-In XOR~
219 491 113 0 3 22
0 18 11 9
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U8A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
5616 0 0
2
5.89968e-315 0
0
14 Logic Display~
6 1109 18 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
5.89968e-315 0
0
14 Logic Display~
6 889 141 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
5.89968e-315 0
0
14 Logic Display~
6 932 244 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
5.89968e-315 0
0
14 Logic Display~
6 994 341 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
5.89968e-315 0
0
14 Logic Display~
6 1056 418 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
5.89968e-315 0
0
14 Logic Display~
6 1065 491 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
5.89968e-315 0
0
14 Logic Display~
6 763 639 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
5.89968e-315 0
0
14 Logic Display~
6 391 647 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
5.89968e-315 0
0
9 Inverter~
13 308 661 0 2 22
0 2 21
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U7B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 7 0
1 U
7100 0 0
2
5.89968e-315 0
0
9 Inverter~
13 600 651 0 2 22
0 13 20
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U7A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 7 0
1 U
3820 0 0
2
5.89968e-315 0
0
9 2-In XOR~
219 589 515 0 3 22
0 13 13 14
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
7678 0 0
2
5.89968e-315 0
0
10 2-In XNOR~
219 587 433 0 3 22
0 13 13 7
0
0 0 624 0
4 4077
-7 -24 21 -16
3 U5A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
961 0 0
2
5.89968e-315 0
0
8 2-In OR~
219 579 157 0 3 22
0 2 13 15
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3178 0 0
2
5.89968e-315 0
0
9 2-In NOR~
219 584 351 0 3 22
0 2 13 19
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3409 0 0
2
5.89968e-315 0
0
10 2-In NAND~
219 591 255 0 3 22
0 2 13 17
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3951 0 0
2
5.89968e-315 0
0
9 2-In AND~
219 584 67 0 3 22
0 2 13 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8885 0 0
2
5.89968e-315 0
0
47
0 1 2 0 0 8320 0 0 18 26 0 4
30 406
30 44
1109 44
1109 36
3 1 3 0 0 4224 0 10 15 0 0 4
488 303
749 303
749 466
757 466
1 3 4 0 0 8320 0 4 12 0 0 3
1084 200
1084 198
1032 198
0 1 5 0 0 8320 0 0 3 0 0 4
810 475
810 293
1085 293
1085 285
0 2 6 0 0 4096 0 0 11 11 0 3
680 691
680 580
742 580
0 1 7 0 0 4096 0 0 11 31 0 3
697 433
697 562
742 562
3 1 8 0 0 4224 0 9 5 0 0 5
685 114
816 114
816 134
876 134
876 99
0 2 2 0 0 0 0 0 9 27 0 3
622 67
622 123
630 123
3 1 9 0 0 4224 0 17 9 0 0 4
524 113
622 113
622 105
630 105
3 1 10 0 0 4224 0 11 6 0 0 3
787 571
1038 571
1038 568
3 1 6 0 0 4224 0 8 7 0 0 3
520 691
946 691
946 635
0 1 11 0 0 4096 0 0 10 22 0 4
301 207
425 207
425 294
433 294
2 2 12 0 0 8320 0 8 10 0 0 4
465 700
425 700
425 312
433 312
0 1 13 0 0 8192 0 0 8 35 0 3
145 570
145 682
465 682
2 0 14 0 0 4096 0 15 0 0 32 3
757 484
656 484
656 515
0 1 15 0 0 8192 0 0 12 28 0 3
849 157
849 189
987 189
3 2 16 0 0 4224 0 16 12 0 0 4
780 205
979 205
979 207
987 207
2 0 17 0 0 4096 0 16 0 0 29 3
731 214
643 214
643 255
1 0 15 0 0 0 0 16 0 0 28 3
731 196
656 196
656 157
1 0 2 0 0 0 0 13 0 0 24 2
248 198
153 198
2 0 13 0 0 0 0 13 0 0 42 3
248 216
244 216
244 264
2 3 11 0 0 4224 0 17 13 0 0 4
475 122
301 122
301 207
293 207
3 1 18 0 0 4224 0 14 17 0 0 4
220 111
467 111
467 104
475 104
0 2 2 0 0 0 0 0 14 43 0 3
153 246
153 120
175 120
1 0 13 0 0 0 0 14 0 0 46 2
175 102
100 102
0 1 2 0 0 0 0 0 26 47 0 4
84 406
30 406
30 661
293 661
3 1 2 0 0 128 0 33 18 0 0 3
605 67
1109 67
1109 36
3 1 15 0 0 4224 0 30 19 0 0 5
612 157
877 157
877 167
889 167
889 159
3 1 17 0 0 4224 0 32 20 0 0 5
618 255
920 255
920 270
932 270
932 262
3 1 19 0 0 4224 0 31 21 0 0 5
623 351
982 351
982 367
994 367
994 359
3 1 7 0 0 4224 0 29 22 0 0 5
626 433
1044 433
1044 444
1056 444
1056 436
3 1 14 0 0 4224 0 28 23 0 0 3
622 515
1065 515
1065 509
2 1 20 0 0 4224 0 27 24 0 0 5
621 651
751 651
751 665
763 665
763 657
2 1 21 0 0 4224 0 26 25 0 0 5
329 661
379 661
379 673
391 673
391 665
0 1 13 0 0 4096 0 0 27 46 0 4
100 570
577 570
577 651
585 651
2 0 13 0 0 0 0 28 0 0 46 2
573 524
100 524
1 0 13 0 0 0 0 28 0 0 46 2
573 506
100 506
2 0 13 0 0 0 0 29 0 0 46 4
571 442
105 442
105 443
100 443
1 0 13 0 0 0 0 29 0 0 46 2
571 424
100 424
2 0 13 0 0 0 0 31 0 0 46 2
571 360
100 360
1 0 2 0 0 128 0 31 0 0 47 2
571 342
84 342
2 0 13 0 0 0 0 32 0 0 46 2
567 264
100 264
1 0 2 0 0 0 0 32 0 0 47 2
567 246
84 246
2 0 13 0 0 0 0 30 0 0 46 2
566 166
100 166
1 0 2 0 0 0 0 30 0 0 47 2
566 148
84 148
1 2 13 0 0 8320 0 2 33 0 0 4
81 585
100 585
100 76
560 76
1 1 2 0 0 0 0 1 33 0 0 3
84 512
84 58
560 58
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
320 26 405 50
330 34 394 50
8 AND Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
314 117 391 141
324 125 380 141
7 OR Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
311 214 404 238
321 222 393 238
9 NAND Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
313 306 398 330
323 314 387 330
8 NOR Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
306 390 399 414
316 398 388 414
9 XNOR Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
306 473 391 497
316 481 380 497
8 XOR Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
159 610 244 634
169 618 233 634
8 NOT Gate
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
