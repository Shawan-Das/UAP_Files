CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
1100 750 1 110 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
72
13 Logic Switch~
5 2026 1029 0 1 11
0 3
0
0 0 21360 180
2 0V
-7 -16 7 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9196 0 0
2
44301.5 1
0
13 Logic Switch~
5 2028 1117 0 1 11
0 2
0
0 0 21360 180
2 0V
-7 -16 7 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3857 0 0
2
44301.5 0
0
13 Logic Switch~
5 1746 1180 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-8 16 6 24
3 D14
-32 7 -11 15
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7125 0 0
2
44301.5 11
0
13 Logic Switch~
5 1880 1195 0 1 11
0 7
0
0 0 21360 90
2 0V
11 0 25 8
3 D13
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3641 0 0
2
44301.5 10
0
13 Logic Switch~
5 1642 1203 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
3 D10
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9821 0 0
2
44301.5 4
0
13 Logic Switch~
5 1507 1201 0 1 11
0 14
0
0 0 21360 90
2 0V
11 0 25 8
2 D9
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3187 0 0
2
44301.5 3
0
13 Logic Switch~
5 1378 1200 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 D8
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
762 0 0
2
44301.5 2
0
13 Logic Switch~
5 1244 1185 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-8 16 6 24
2 D7
-29 7 -15 15
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
39 0 0
2
44301.5 1
0
13 Logic Switch~
5 295 564 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-32 0 -18 8
1 D
-27 -10 -20 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9450 0 0
2
44301.5 0
0
13 Logic Switch~
5 851 556 0 1 11
0 22
0
0 0 21360 180
2 0V
-7 -16 7 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3236 0 0
2
44301.5 1
0
13 Logic Switch~
5 853 644 0 1 11
0 21
0
0 0 21360 180
2 0V
-7 -16 7 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3321 0 0
2
44301.5 2
0
13 Logic Switch~
5 1113 662 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8879 0 0
2
44301.5 3
0
13 Logic Switch~
5 1691 295 0 1 11
0 27
0
0 0 21360 180
2 0V
-7 -16 7 -8
2 V8
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5433 0 0
2
44301.5 4
0
13 Logic Switch~
5 1048 575 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3679 0 0
2
44301.5 5
0
13 Logic Switch~
5 1111 525 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9342 0 0
2
44301.5 6
0
13 Logic Switch~
5 338 326 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-32 0 -18 8
2 V4
-31 -10 -17 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3623 0 0
2
44301.5 7
0
13 Logic Switch~
5 1149 357 0 10 11
0 45 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-8 16 6 24
2 D0
-29 7 -15 15
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3722 0 0
2
44301.5 8
0
13 Logic Switch~
5 1283 372 0 1 11
0 44
0
0 0 21360 90
2 0V
11 0 25 8
2 D6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8993 0 0
2
44301.5 9
0
13 Logic Switch~
5 1412 373 0 10 11
0 43 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 D5
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3723 0 0
2
44301.5 10
0
13 Logic Switch~
5 1547 375 0 1 11
0 42
0
0 0 21360 90
2 0V
11 0 25 8
2 D4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6244 0 0
2
44301.5 11
0
13 Logic Switch~
5 1689 207 0 1 11
0 28
0
0 0 21360 180
2 0V
-7 -16 7 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6421 0 0
2
44301.5 12
0
13 Logic Switch~
5 442 328 0 1 11
0 46
0
0 0 21360 90
2 0V
-5 22 9 30
3 DSL
15 22 36 30
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7743 0 0
2
44301.5 13
0
13 Logic Switch~
5 423 330 0 10 11
0 36 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-10 19 4 27
3 DSR
-41 20 -20 28
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9840 0 0
2
44301.5 14
0
13 Logic Switch~
5 362 189 0 10 11
0 57 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 S1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6910 0 0
2
44301.5 15
0
13 Logic Switch~
5 398 187 0 1 11
0 56
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 S0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
449 0 0
2
44301.5 16
0
13 Logic Switch~
5 664 155 0 1 11
0 48
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 D0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8761 0 0
2
44301.5 17
0
13 Logic Switch~
5 628 155 0 10 11
0 49 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 D1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6748 0 0
2
44301.5 18
0
13 Logic Switch~
5 600 156 0 1 11
0 50
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 D2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7393 0 0
2
44301.5 19
0
13 Logic Switch~
5 568 154 0 10 11
0 51 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 D3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7699 0 0
2
44301.5 20
0
14 Logic Display~
6 1614 930 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6638 0 0
2
44301.5 5
0
14 Logic Display~
6 1579 930 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L18
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4595 0 0
2
44301.5 4
0
5 4013~
219 1938 1108 0 6 22
0 3 7 4 2 58 5
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U10B
19 -61 47 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 9 0
1 U
9395 0 0
2
44301.5 1
0
5 4013~
219 1800 1111 0 6 22
0 3 8 4 2 59 6
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U10A
19 -61 47 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 9 0
1 U
3303 0 0
2
44301.5 0
0
5 4013~
219 1294 1114 0 6 22
0 3 16 4 2 60 12
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U9B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 8 0
1 U
4498 0 0
2
44301.5 14
0
5 4013~
219 1436 1113 0 6 22
0 3 15 4 2 61 11
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U9A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 8 0
1 U
9728 0 0
2
44301.5 13
0
5 4013~
219 1572 1113 0 6 22
0 3 14 4 2 62 10
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U8B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 7 0
1 U
3789 0 0
2
44301.5 12
0
5 4013~
219 1698 1107 0 6 22
0 3 13 4 2 63 9
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U8A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 7 0
1 U
3978 0 0
2
44301.5 11
0
7 Pulser~
4 1165 1090 0 10 12
0 4 64 4 65 0 0 5 5 1
8
0
0 0 4656 0
0
3 V15
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3494 0 0
2
44301.5 10
0
14 Logic Display~
6 1471 933 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3507 0 0
2
44301.5 9
0
14 Logic Display~
6 1495 933 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5151 0 0
2
44301.5 8
0
14 Logic Display~
6 1519 934 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3701 0 0
2
44301.5 7
0
14 Logic Display~
6 1547 933 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8585 0 0
2
44301.5 6
0
5 4013~
219 361 635 0 6 22
0 22 17 24 21 66 20
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U7B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 6 0
1 U
8809 0 0
2
44301.5 21
0
5 4013~
219 503 634 0 6 22
0 22 20 24 21 67 19
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U7A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 6 0
1 U
5993 0 0
2
44301.5 22
0
5 4013~
219 639 634 0 6 22
0 22 19 24 21 68 18
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U6B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 5 0
1 U
8654 0 0
2
44301.5 23
0
5 4013~
219 769 631 0 6 22
0 22 18 24 21 69 23
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U6A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 5 0
1 U
7223 0 0
2
44301.5 24
0
7 Pulser~
4 232 611 0 10 12
0 24 70 24 71 0 0 5 5 1
8
0
0 0 4656 0
0
3 V12
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3641 0 0
2
44301.5 25
0
14 Logic Display~
6 538 454 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3104 0 0
2
44301.5 26
0
14 Logic Display~
6 562 454 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3296 0 0
2
44301.5 27
0
14 Logic Display~
6 586 455 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8534 0 0
2
44301.5 28
0
14 Logic Display~
6 614 454 0 1 2
10 23
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
949 0 0
2
44301.5 29
0
14 Logic Display~
6 1640 493 0 1 2
10 29
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3371 0 0
2
44301.5 30
0
5 4013~
219 1167 611 0 6 22
0 26 30 34 25 72 33
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U5B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 4 0
1 U
7311 0 0
2
44301.5 31
0
5 4013~
219 1309 611 0 6 22
0 26 33 34 25 73 32
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U5A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 4 0
1 U
3409 0 0
2
44301.5 32
0
5 4013~
219 1445 611 0 6 22
0 26 32 34 25 74 31
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U4B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 3 0
1 U
3526 0 0
2
44301.5 33
0
5 4013~
219 1575 611 0 6 22
0 26 31 34 25 75 29
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U4A
15 -64 36 -56
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 3 0
1 U
4129 0 0
2
44301.5 34
0
7 Pulser~
4 1042 632 0 10 12
0 34 76 34 77 0 0 5 5 1
8
0
0 0 4656 0
0
2 V6
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6278 0 0
2
44301.5 35
0
14 Logic Display~
6 1452 105 0 1 2
10 37
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3482 0 0
2
44301.5 36
0
14 Logic Display~
6 1424 106 0 1 2
10 38
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8323 0 0
2
44301.5 37
0
14 Logic Display~
6 1400 105 0 1 2
10 39
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3984 0 0
2
44301.5 38
0
14 Logic Display~
6 1376 105 0 1 2
10 40
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7622 0 0
2
44301.5 39
0
7 Pulser~
4 1070 262 0 10 12
0 41 78 41 79 0 0 5 5 1
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
816 0 0
2
44301.5 40
0
5 4013~
219 1607 282 0 6 22
0 28 42 41 27 80 37
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U3B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 2 0
1 U
4656 0 0
2
44301.5 41
0
5 4013~
219 1477 285 0 6 22
0 28 43 41 27 81 38
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U3A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 2 0
1 U
6356 0 0
2
44301.5 42
0
5 4013~
219 1341 285 0 6 22
0 28 44 41 27 82 39
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U2B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 1 0
1 U
7479 0 0
2
44301.5 43
0
5 4013~
219 1199 286 0 6 22
0 28 45 41 27 83 40
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U2A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 1 0
1 U
5690 0 0
2
44301.5 44
0
7 74LS194
49 510 249 0 14 29
0 47 57 56 36 46 35 51 50 49
48 52 53 54 55
0
0 0 4848 0
6 74F194
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 10 9 2 7 1 6 5 4
3 12 13 14 15 11 10 9 2 7
1 6 5 4 3 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
5617 0 0
2
44301.5 45
0
14 Logic Display~
6 692 206 0 1 2
10 52
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3903 0 0
2
44301.5 46
0
14 Logic Display~
6 716 206 0 1 2
10 53
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4452 0 0
2
44301.5 47
0
14 Logic Display~
6 740 207 0 1 2
10 54
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6282 0 0
2
44301.5 48
0
14 Logic Display~
6 768 206 0 1 2
10 55
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7187 0 0
2
44301.5 49
0
7 Pulser~
4 371 294 0 10 12
0 47 84 47 85 0 0 5 5 1
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6866 0 0
2
44301.5 50
0
107
1 0 2 0 0 4096 0 2 0 0 6 4
2014 1117
1972 1117
1972 1125
1938 1125
0 1 3 0 0 8192 0 0 1 4 0 3
1938 1026
1938 1029
2012 1029
1 0 3 0 0 0 0 33 0 0 4 2
1800 1054
1800 1026
0 0 3 0 0 4096 0 0 0 32 13 2
1698 1026
1938 1026
4 0 2 0 0 0 0 33 0 0 6 2
1800 1117
1800 1141
0 4 2 0 0 4096 0 0 32 29 0 3
1698 1141
1938 1141
1938 1114
3 0 4 0 0 8192 0 33 0 0 8 3
1776 1093
1772 1093
1772 1122
0 3 4 0 0 8192 0 0 32 21 0 5
1670 1125
1670 1122
1906 1122
1906 1090
1914 1090
6 1 5 0 0 8320 0 32 30 0 0 4
1962 1072
1962 961
1614 961
1614 948
6 1 6 0 0 12416 0 33 31 0 0 5
1824 1075
1845 1075
1845 966
1579 966
1579 948
1 2 7 0 0 4224 0 4 32 0 0 3
1881 1182
1881 1072
1914 1072
1 2 8 0 0 4224 0 3 33 0 0 3
1747 1167
1747 1075
1776 1075
1 0 3 0 0 0 0 32 0 0 0 2
1938 1051
1938 1020
6 1 9 0 0 12416 0 37 42 0 0 5
1722 1071
1736 1071
1736 977
1547 977
1547 951
6 1 10 0 0 12416 0 36 41 0 0 5
1596 1077
1606 1077
1606 993
1519 993
1519 952
6 1 11 0 0 8320 0 35 40 0 0 3
1460 1077
1495 1077
1495 951
6 1 12 0 0 12416 0 34 39 0 0 5
1318 1078
1343 1078
1343 986
1471 986
1471 951
3 0 4 0 0 0 0 36 0 0 21 3
1548 1095
1545 1095
1545 1125
3 0 4 0 0 0 0 35 0 0 21 3
1412 1095
1408 1095
1408 1125
3 0 4 0 0 0 0 34 0 0 21 3
1270 1096
1266 1096
1266 1125
0 3 4 0 0 12416 0 0 37 22 0 6
1203 1080
1222 1080
1222 1125
1670 1125
1670 1089
1674 1089
1 3 4 0 0 0 0 38 38 0 0 6
1141 1081
1131 1081
1131 1067
1203 1067
1203 1081
1189 1081
1 2 13 0 0 8320 0 5 37 0 0 4
1643 1190
1644 1190
1644 1071
1674 1071
1 2 14 0 0 4224 0 6 36 0 0 3
1508 1188
1508 1077
1548 1077
1 2 15 0 0 4224 0 7 35 0 0 3
1379 1187
1379 1077
1412 1077
1 2 16 0 0 4224 0 8 34 0 0 3
1245 1172
1245 1078
1270 1078
1 0 3 0 0 0 0 35 0 0 32 2
1436 1056
1436 1025
1 0 3 0 0 0 0 36 0 0 32 2
1572 1056
1572 1025
4 4 2 0 0 8320 0 37 34 0 0 4
1698 1113
1698 1143
1294 1143
1294 1120
4 0 2 0 0 0 0 36 0 0 29 2
1572 1119
1572 1143
4 0 2 0 0 0 0 35 0 0 29 2
1436 1119
1436 1143
1 1 3 0 0 8320 0 37 34 0 0 4
1698 1050
1698 1025
1294 1025
1294 1057
1 2 17 0 0 8320 0 9 43 0 0 4
307 564
329 564
329 599
337 599
0 2 18 0 0 8192 0 0 46 40 0 3
673 598
673 595
745 595
0 2 19 0 0 4096 0 0 45 41 0 2
562 598
615 598
0 2 20 0 0 8192 0 0 44 42 0 3
410 599
410 598
479 598
1 0 21 0 0 4096 0 11 0 0 50 2
839 644
769 644
1 0 22 0 0 4096 0 10 0 0 53 2
837 556
769 556
6 1 23 0 0 12416 0 46 51 0 0 5
793 595
803 595
803 498
614 498
614 472
6 1 18 0 0 12416 0 45 50 0 0 5
663 598
673 598
673 514
586 514
586 473
6 1 19 0 0 8320 0 44 49 0 0 3
527 598
562 598
562 472
6 1 20 0 0 12416 0 43 48 0 0 5
385 599
410 599
410 507
538 507
538 472
3 0 24 0 0 8192 0 45 0 0 46 3
615 616
612 616
612 646
3 0 24 0 0 0 0 44 0 0 46 3
479 616
475 616
475 646
3 0 24 0 0 0 0 43 0 0 46 3
337 617
333 617
333 646
0 3 24 0 0 12416 0 0 46 47 0 6
270 601
289 601
289 646
737 646
737 613
745 613
1 3 24 0 0 0 0 47 47 0 0 6
208 602
198 602
198 588
270 588
270 602
256 602
1 0 22 0 0 0 0 44 0 0 53 2
503 577
503 546
1 0 22 0 0 0 0 45 0 0 53 2
639 577
639 546
4 4 21 0 0 8320 0 46 43 0 0 4
769 637
769 664
361 664
361 641
4 0 21 0 0 0 0 45 0 0 50 2
639 640
639 664
4 0 21 0 0 0 0 44 0 0 50 2
503 640
503 664
1 1 22 0 0 8320 0 46 43 0 0 4
769 574
769 546
361 546
361 578
1 0 25 0 0 4096 0 12 0 0 70 3
1125 662
1168 662
1168 641
1 0 26 0 0 4096 0 53 0 0 73 2
1167 554
1167 525
1 0 27 0 0 4096 0 13 0 0 91 2
1677 295
1607 295
1 0 28 0 0 4096 0 21 0 0 94 2
1675 207
1607 207
6 1 29 0 0 8320 0 56 52 0 0 3
1599 575
1640 575
1640 511
1 2 30 0 0 4224 0 14 53 0 0 2
1060 575
1143 575
6 2 31 0 0 4224 0 55 56 0 0 2
1469 575
1551 575
6 2 32 0 0 4224 0 54 55 0 0 2
1333 575
1421 575
6 2 33 0 0 4224 0 53 54 0 0 2
1191 575
1285 575
3 0 34 0 0 8192 0 55 0 0 66 3
1421 593
1418 593
1418 622
3 0 34 0 0 0 0 54 0 0 66 3
1285 593
1281 593
1281 622
3 0 34 0 0 0 0 53 0 0 66 3
1143 593
1139 593
1139 622
0 3 34 0 0 12416 0 0 56 67 0 6
1076 623
1095 623
1095 622
1543 622
1543 593
1551 593
1 3 34 0 0 0 0 57 57 0 0 6
1018 623
1004 623
1004 597
1076 597
1076 623
1066 623
1 0 26 0 0 0 0 54 0 0 73 2
1309 554
1309 525
1 0 26 0 0 0 0 55 0 0 73 2
1445 554
1445 525
4 4 25 0 0 8320 0 56 53 0 0 4
1575 617
1575 641
1167 641
1167 617
4 0 25 0 0 0 0 55 0 0 70 2
1445 617
1445 641
4 0 25 0 0 0 0 54 0 0 70 2
1309 617
1309 641
1 1 26 0 0 8320 0 56 15 0 0 3
1575 554
1575 525
1123 525
1 6 35 0 0 8320 0 16 67 0 0 5
350 326
350 325
414 325
414 285
472 285
1 4 36 0 0 4224 0 23 67 0 0 3
424 317
424 258
478 258
6 1 37 0 0 12416 0 63 58 0 0 5
1631 246
1641 246
1641 149
1452 149
1452 123
6 1 38 0 0 12416 0 64 59 0 0 5
1501 249
1511 249
1511 165
1424 165
1424 124
6 1 39 0 0 8320 0 65 60 0 0 3
1365 249
1400 249
1400 123
6 1 40 0 0 12416 0 66 61 0 0 5
1223 250
1248 250
1248 158
1376 158
1376 123
3 0 41 0 0 8192 0 64 0 0 83 3
1453 267
1450 267
1450 297
3 0 41 0 0 0 0 65 0 0 83 3
1317 267
1313 267
1313 297
3 0 41 0 0 0 0 66 0 0 83 3
1175 268
1171 268
1171 297
0 3 41 0 0 12416 0 0 63 84 0 6
1108 252
1127 252
1127 297
1575 297
1575 264
1583 264
1 3 41 0 0 0 0 62 62 0 0 6
1046 253
1036 253
1036 239
1108 239
1108 253
1094 253
1 2 42 0 0 8320 0 20 63 0 0 4
1548 362
1549 362
1549 246
1583 246
1 2 43 0 0 4224 0 19 64 0 0 3
1413 360
1413 249
1453 249
1 2 44 0 0 4224 0 18 65 0 0 3
1284 359
1284 249
1317 249
1 2 45 0 0 4224 0 17 66 0 0 3
1150 344
1150 250
1175 250
1 0 28 0 0 0 0 65 0 0 94 2
1341 228
1341 197
1 0 28 0 0 0 0 64 0 0 94 2
1477 228
1477 197
4 4 27 0 0 8320 0 63 66 0 0 4
1607 288
1607 315
1199 315
1199 292
4 0 27 0 0 0 0 64 0 0 91 2
1477 291
1477 315
4 0 27 0 0 0 0 65 0 0 91 2
1341 291
1341 315
1 1 28 0 0 8320 0 63 66 0 0 4
1607 225
1607 197
1199 197
1199 229
1 5 46 0 0 4224 0 22 67 0 0 3
443 315
443 267
478 267
0 1 47 0 0 8320 0 0 67 97 0 4
396 278
416 278
416 213
478 213
1 3 47 0 0 0 0 72 72 0 0 6
347 285
342 285
342 271
396 271
396 285
395 285
1 10 48 0 0 8320 0 26 67 0 0 3
664 167
664 240
542 240
1 9 49 0 0 8320 0 27 67 0 0 3
628 167
628 231
542 231
1 8 50 0 0 8320 0 28 67 0 0 3
600 168
600 222
542 222
1 7 51 0 0 4224 0 29 67 0 0 3
568 166
568 213
542 213
11 1 52 0 0 4224 0 67 68 0 0 3
542 258
692 258
692 224
12 1 53 0 0 4224 0 67 69 0 0 3
542 267
716 267
716 224
13 1 54 0 0 4224 0 67 70 0 0 3
542 276
740 276
740 225
14 1 55 0 0 4224 0 67 71 0 0 3
542 285
768 285
768 224
1 3 56 0 0 8320 0 25 67 0 0 3
398 199
398 240
478 240
1 2 57 0 0 8320 0 24 67 0 0 3
362 201
362 231
478 231
15
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
1576 1235 1629 1263
1584 1242 1620 1260
4 PIPO
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
185 211 250 237
194 219 240 237
5 DSP=1
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
186 238 251 264
195 245 241 263
5 DSL=1
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
119 238 176 264
129 245 165 263
4 LEST
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
121 210 186 236
130 218 176 236
5 RIGHT
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
38 179 111 205
47 186 101 204
6 0    0
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
37 211 110 237
46 218 100 236
6 0    1
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
40 238 113 264
49 246 103 264
6 1    0
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
40 265 113 291
49 272 103 290
6 1    1
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 7
30 139 114 165
40 147 103 165
7 S1   S0
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
527 682 580 710
535 688 571 706
4 SIPO
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
1336 660 1389 688
1344 667 1380 685
4 SISO
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
1345 401 1398 429
1353 408 1389 426
4 PIPO
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 15
496 304 646 332
503 309 638 327
15 Universal Shift
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 8
650 300 743 328
660 308 732 326
8 Resister
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
