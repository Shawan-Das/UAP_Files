CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 237 408 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-8 16 6 24
2 D7
-6 30 8 38
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7670 0 0
2
44301.5 7
0
13 Logic Switch~
5 371 423 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-8 14 6 22
2 D8
-8 24 6 32
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
951 0 0
2
44301.5 6
0
13 Logic Switch~
5 500 424 0 1 11
0 14
0
0 0 21360 90
2 0V
-5 13 9 21
2 D9
-3 27 11 35
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9536 0 0
2
44301.5 5
0
13 Logic Switch~
5 635 426 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-7 15 7 23
3 D10
-4 29 17 37
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5495 0 0
2
44301.5 4
0
13 Logic Switch~
5 873 418 0 1 11
0 7
0
0 0 21360 90
2 0V
-4 15 10 23
3 D13
-7 28 14 36
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8152 0 0
2
44301.5 3
0
13 Logic Switch~
5 739 403 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-8 16 6 24
3 D14
-10 34 11 42
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6223 0 0
2
44301.5 2
0
13 Logic Switch~
5 1021 340 0 1 11
0 2
0
0 0 21360 180
2 0V
-7 -16 7 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5441 0 0
2
44301.5 1
0
13 Logic Switch~
5 1019 252 0 1 11
0 3
0
0 0 21360 180
2 0V
-7 -16 7 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3189 0 0
2
44301.5 0
0
14 Logic Display~
6 540 156 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8460 0 0
2
44301.5 20
0
14 Logic Display~
6 512 157 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5179 0 0
2
44301.5 19
0
14 Logic Display~
6 488 156 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3593 0 0
2
44301.5 18
0
14 Logic Display~
6 464 156 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3928 0 0
2
44301.5 17
0
7 Pulser~
4 158 313 0 10 12
0 4 17 4 18 0 0 5 5 5
8
0
0 0 4656 0
0
3 V15
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
363 0 0
2
44301.5 16
0
5 4013~
219 691 330 0 6 22
0 3 13 4 2 19 9
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U3B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 3 0
1 U
8132 0 0
2
44301.5 15
0
5 4013~
219 565 336 0 6 22
0 3 14 4 2 20 10
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U3A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 3 0
1 U
65 0 0
2
44301.5 14
0
5 4013~
219 429 336 0 6 22
0 3 15 4 2 21 11
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U2B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 2 0
1 U
6609 0 0
2
44301.5 13
0
5 4013~
219 287 337 0 6 22
0 3 16 4 2 22 12
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U2A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 2 0
1 U
8995 0 0
2
44301.5 12
0
5 4013~
219 793 334 0 6 22
0 3 8 4 2 23 6
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 1 0
1 U
3918 0 0
2
44301.5 11
0
5 4013~
219 931 331 0 6 22
0 3 7 4 2 24 5
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 1 0
1 U
7519 0 0
2
44301.5 10
0
14 Logic Display~
6 572 153 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L18
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
377 0 0
2
44301.5 9
0
14 Logic Display~
6 607 153 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8816 0 0
2
44301.5 8
0
32
1 0 2 0 0 4096 0 7 0 0 6 4
1007 340
965 340
965 348
931 348
0 1 3 0 0 8192 0 0 8 4 0 3
931 249
931 252
1005 252
1 0 3 0 0 0 0 18 0 0 4 2
793 277
793 249
0 0 3 0 0 4096 0 0 0 32 13 2
691 249
931 249
4 0 2 0 0 0 0 18 0 0 6 2
793 340
793 364
0 4 2 0 0 4096 0 0 19 29 0 3
691 364
931 364
931 337
3 0 4 0 0 8192 0 18 0 0 8 3
769 316
765 316
765 345
0 3 4 0 0 8192 0 0 19 21 0 5
663 348
663 345
899 345
899 313
907 313
6 1 5 0 0 8336 0 19 21 0 0 4
955 295
955 181
607 181
607 171
6 1 6 0 0 12416 0 18 20 0 0 5
817 298
838 298
838 189
572 189
572 171
1 2 7 0 0 4224 0 5 19 0 0 3
874 405
874 295
907 295
1 2 8 0 0 4224 0 6 18 0 0 3
740 390
740 298
769 298
1 0 3 0 0 0 0 19 0 0 0 2
931 274
931 243
6 1 9 0 0 12416 0 14 9 0 0 5
715 294
729 294
729 200
540 200
540 174
6 1 10 0 0 12416 0 15 10 0 0 5
589 300
599 300
599 216
512 216
512 175
6 1 11 0 0 8320 0 16 11 0 0 3
453 300
488 300
488 174
6 1 12 0 0 12416 0 17 12 0 0 5
311 301
336 301
336 209
464 209
464 174
3 0 4 0 0 0 0 15 0 0 21 3
541 318
538 318
538 348
3 0 4 0 0 0 0 16 0 0 21 3
405 318
401 318
401 348
3 0 4 0 0 0 0 17 0 0 21 3
263 319
259 319
259 348
0 3 4 0 0 12416 0 0 14 22 0 6
196 303
215 303
215 348
663 348
663 312
667 312
1 3 4 0 0 0 0 13 13 0 0 6
134 304
124 304
124 290
196 290
196 304
182 304
1 2 13 0 0 8320 0 4 14 0 0 4
636 413
637 413
637 294
667 294
1 2 14 0 0 4224 0 3 15 0 0 3
501 411
501 300
541 300
1 2 15 0 0 4224 0 2 16 0 0 3
372 410
372 300
405 300
1 2 16 0 0 4224 0 1 17 0 0 3
238 395
238 301
263 301
1 0 3 0 0 0 0 16 0 0 32 2
429 279
429 248
1 0 3 0 0 0 0 15 0 0 32 2
565 279
565 248
4 4 2 0 0 8320 0 14 17 0 0 4
691 336
691 366
287 366
287 343
4 0 2 0 0 0 0 15 0 0 29 2
565 342
565 366
4 0 2 0 0 0 0 16 0 0 29 2
429 342
429 366
1 1 3 0 0 8320 0 14 17 0 0 4
691 273
691 248
287 248
287 280
1
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
569 458 622 486
577 465 613 483
4 PIPO
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
