CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
20
13 Logic Switch~
5 175 40 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89969e-315 0
0
13 Logic Switch~
5 106 39 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
99 -138 113 -130
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89969e-315 0
0
13 Logic Switch~
5 29 41 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89969e-315 0
0
5 7415~
219 462 237 0 4 22
0 2 3 5 6
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 6 0
1 U
3421 0 0
2
5.89969e-315 0
0
8 4-In OR~
219 592 173 0 5 22
0 12 13 11 6 4
0
0 0 608 0
4 4072
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
8157 0 0
2
5.89969e-315 0
0
9 2-In AND~
219 458 372 0 3 22
0 2 5 8
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
5572 0 0
2
5.89969e-315 0
0
9 2-In AND~
219 460 330 0 3 22
0 3 5 10
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
8901 0 0
2
5.89969e-315 0
0
9 2-In AND~
219 461 291 0 3 22
0 2 3 9
0
0 0 608 0
5 74F08
-18 -24 17 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
7361 0 0
2
5.89969e-315 0
0
8 3-In OR~
219 597 330 0 4 22
0 9 10 8 7
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U2B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 2 0
1 U
4747 0 0
2
5.89969e-315 5.26354e-315
0
14 Logic Display~
6 673 326 0 1 2
10 7
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L5
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
5.89969e-315 0
0
14 Logic Display~
6 665 169 0 1 2
10 4
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L4
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
5.89969e-315 0
0
9 Inverter~
13 229 200 0 2 22
0 5 14
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
9998 0 0
2
5.89969e-315 0
0
9 Inverter~
13 150 154 0 2 22
0 3 15
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
3536 0 0
2
5.89969e-315 0
0
9 Inverter~
13 71 105 0 2 22
0 2 16
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
4597 0 0
2
5.89969e-315 0
0
5 7415~
219 458 191 0 4 22
0 2 3 14 11
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 1 0
1 U
3835 0 0
2
5.89969e-315 0
0
5 7415~
219 457 154 0 4 22
0 2 15 5 13
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 1 0
1 U
3670 0 0
2
5.89969e-315 0
0
5 7415~
219 459 114 0 4 22
0 16 3 5 12
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 1 0
1 U
5616 0 0
2
5.89969e-315 0
0
14 Logic Display~
6 194 440 0 1 2
10 5
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L3
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
5.89969e-315 0
0
14 Logic Display~
6 117 441 0 1 2
10 3
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L2
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
5.89969e-315 0
0
14 Logic Display~
6 40 441 0 1 2
10 2
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
5.89969e-315 0
0
33
1 0 2 0 0 4096 0 15 0 0 33 2
434 182
40 182
2 0 3 0 0 4096 0 15 0 0 32 2
434 191
117 191
5 1 4 0 0 4224 0 5 11 0 0 2
625 173
649 173
1 0 2 0 0 0 0 16 0 0 33 2
433 145
40 145
3 0 5 0 0 4096 0 4 0 0 31 2
438 246
194 246
2 0 3 0 0 4096 0 4 0 0 32 2
438 237
117 237
1 0 2 0 0 4096 0 4 0 0 33 2
438 228
40 228
4 4 6 0 0 8320 0 4 5 0 0 5
483 237
483 200
551 200
551 187
575 187
2 0 5 0 0 0 0 6 0 0 31 2
434 381
194 381
1 0 2 0 0 0 0 6 0 0 33 2
434 363
40 363
2 0 5 0 0 0 0 7 0 0 31 2
436 339
194 339
1 0 3 0 0 0 0 7 0 0 32 2
436 321
117 321
2 0 3 0 0 0 0 8 0 0 32 2
437 300
117 300
1 0 2 0 0 0 0 8 0 0 33 2
437 282
40 282
1 4 7 0 0 4224 0 10 9 0 0 2
657 330
630 330
3 3 8 0 0 4224 0 6 9 0 0 4
479 372
556 372
556 339
584 339
3 1 9 0 0 4224 0 8 9 0 0 4
482 291
556 291
556 321
584 321
3 2 10 0 0 4224 0 7 9 0 0 2
481 330
585 330
3 0 5 0 0 0 0 16 0 0 31 2
433 163
194 163
3 0 5 0 0 0 0 17 0 0 31 2
435 123
194 123
2 0 3 0 0 0 0 17 0 0 32 2
435 114
117 114
4 3 11 0 0 4224 0 15 5 0 0 4
479 191
540 191
540 178
575 178
4 1 12 0 0 12416 0 17 5 0 0 6
480 114
484 114
484 146
550 146
550 160
575 160
4 2 13 0 0 4224 0 16 5 0 0 4
478 154
541 154
541 169
575 169
2 3 14 0 0 4224 0 12 15 0 0 2
250 200
434 200
1 0 5 0 0 0 0 12 0 0 31 2
214 200
194 200
2 2 15 0 0 4224 0 13 16 0 0 2
171 154
433 154
1 0 3 0 0 0 0 13 0 0 32 2
135 154
117 154
2 1 16 0 0 4224 0 14 17 0 0 2
92 105
435 105
1 0 2 0 0 0 0 14 0 0 33 2
56 105
40 105
1 1 5 0 0 8320 0 1 18 0 0 3
187 40
194 40
194 426
1 1 3 0 0 8336 0 2 19 0 0 3
118 39
117 39
117 427
1 1 2 0 0 8320 0 3 20 0 0 3
41 41
40 41
40 427
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
