CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
320 0 25 150 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.326954 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 85 303 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 1 0 -1 0
1 V
961 0 0
2
5.89975e-315 0
0
9 2-In AND~
219 1064 360 0 3 22
0 7 8 9
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U5B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3178 0 0
2
44256.4 0
0
8 2-In OR~
219 920 335 0 3 22
0 11 9 10
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3409 0 0
2
44256.4 0
0
9 2-In AND~
219 829 263 0 3 22
0 4 3 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3951 0 0
2
44256.4 0
0
12 Hex Display~
7 951 62 0 18 19
10 6 4 5 21 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP4
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
8885 0 0
2
44256.4 4
0
7 74LS293
154 955 219 0 8 17
0 11 11 22 7 5 4 6 23
0
0 0 4848 90
7 74LS293
-24 -35 25 -27
2 U4
248 -146 262 -138
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 512 1 0 0 0
1 U
3780 0 0
2
44256.4 3
0
7 74LS293
154 1008 219 0 8 17
0 10 10 2 12 7 3 8 12
0
0 0 4848 90
7 74LS293
-24 -35 25 -27
2 U3
203 -124 217 -116
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 0 1 0 0 0
1 U
9265 0 0
2
44256.4 2
0
12 Hex Display~
7 984 62 0 18 19
10 12 8 3 7 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9442 0 0
2
44256.4 1
0
7 Pulser~
4 778 351 0 10 12
0 24 25 26 27 0 0 5 5 1
8
0
0 0 4656 0
0
2 V3
-4 -51 10 -43
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9424 0 0
2
44256.4 0
0
7 Pulser~
4 123 248 0 10 12
0 15 28 15 29 0 0 5 5 1
8
0
0 0 4656 0
0
2 V2
-4 -51 10 -43
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9968 0 0
2
5.89975e-315 0
0
12 Hex Display~
7 380 69 0 18 19
10 19 14 16 13 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9281 0 0
2
5.89975e-315 0
0
7 74LS293
154 478 230 0 8 17
0 2 17 30 13 2 17 18 31
0
0 0 4848 0
7 74LS293
-24 -35 25 -27
2 U2
-7 -36 7 -28
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 512 1 0 0 0
1 U
8464 0 0
2
5.89975e-315 0
0
7 74LS293
154 269 230 0 8 17
0 13 14 15 19 13 16 14 19
0
0 0 4848 0
7 74LS293
-24 -35 25 -27
2 U1
-7 -36 7 -28
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 0 1 0 0 0
1 U
7168 0 0
2
5.89975e-315 0
0
12 Hex Display~
7 347 69 0 18 19
10 18 17 2 32 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
3171 0 0
2
5.89975e-315 0
0
35
0 3 2 0 0 8320 0 0 7 29 0 4
534 221
534 283
1013 283
1013 255
0 2 3 0 0 4240 0 0 4 18 0 4
981 135
783 135
783 272
805 272
0 1 4 0 0 4224 0 0 4 5 0 4
951 170
797 170
797 254
805 254
5 3 5 0 0 4224 0 6 5 0 0 4
942 185
942 94
948 94
948 86
6 2 4 0 0 0 0 6 5 0 0 4
951 185
951 94
954 94
954 86
7 1 6 0 0 4224 0 6 5 0 0 2
960 185
960 86
0 1 7 0 0 8192 0 0 2 15 0 4
1080 269
1107 269
1107 369
1082 369
0 2 8 0 0 8320 0 0 2 19 0 4
1013 172
1092 172
1092 351
1082 351
2 3 9 0 0 12416 0 3 2 0 0 4
907 344
903 344
903 360
1037 360
0 1 10 0 0 4224 0 0 7 11 0 2
995 335
995 249
3 2 10 0 0 0 0 3 7 0 0 3
953 335
1004 335
1004 249
0 1 11 0 0 4096 0 0 3 14 0 3
883 263
883 326
907 326
1 0 11 0 0 0 0 6 0 0 14 2
942 249
942 263
3 2 11 0 0 4224 0 4 6 0 0 3
850 263
951 263
951 249
0 4 7 0 0 8320 0 0 6 17 0 5
995 156
1080 156
1080 300
969 300
969 255
8 4 12 0 0 12416 0 7 7 0 0 6
1022 185
1022 181
1037 181
1037 263
1022 263
1022 255
4 5 7 0 0 0 0 8 7 0 0 4
975 86
975 156
995 156
995 185
3 6 3 0 0 0 0 8 7 0 0 4
981 86
981 148
1004 148
1004 185
2 7 8 0 0 0 0 8 7 0 0 4
987 86
987 138
1013 138
1013 185
1 8 12 0 0 0 0 8 7 0 0 4
993 86
993 126
1022 126
1022 185
0 4 13 0 0 8192 0 0 12 22 0 4
331 222
331 260
440 260
440 248
0 4 13 0 0 12416 0 0 11 27 0 4
304 221
304 222
371 222
371 93
0 2 14 0 0 8320 0 0 11 24 0 3
314 239
383 239
383 93
2 7 14 0 0 0 0 13 13 0 0 6
237 230
222 230
222 288
314 288
314 239
301 239
3 3 15 0 0 4224 0 10 13 0 0 2
147 239
231 239
1 3 15 0 0 0 0 10 10 0 0 6
99 239
89 239
89 224
161 224
161 239
147 239
5 1 13 0 0 0 0 13 13 0 0 6
301 221
305 221
305 184
223 184
223 221
237 221
6 3 16 0 0 8320 0 13 11 0 0 3
301 230
377 230
377 93
5 3 2 0 0 128 0 12 14 0 0 5
510 221
534 221
534 160
344 160
344 93
6 2 17 0 0 12416 0 12 14 0 0 5
510 230
529 230
529 155
350 155
350 93
7 1 18 0 0 12416 0 12 14 0 0 5
510 239
524 239
524 150
356 150
356 93
0 1 19 0 0 8320 0 0 11 35 0 3
309 248
389 248
389 93
6 2 17 0 0 0 0 12 12 0 0 6
510 230
519 230
519 172
427 172
427 230
446 230
5 1 2 0 0 0 0 12 12 0 0 6
510 221
514 221
514 185
432 185
432 221
446 221
4 8 19 0 0 0 0 13 13 0 0 6
231 248
227 248
227 263
309 263
309 248
301 248
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
