CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
240 460 30 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
59
13 Logic Switch~
5 498 570 0 1 11
0 2
0
0 0 21360 0
2 0V
-31 -4 -17 4
3 C15
-250 -120 -229 -112
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3122 0 0
2
44257.7 0
0
13 Logic Switch~
5 810 904 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-4 27 10 35
2 B1
-5 16 9 24
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6242 0 0
2
44257.6 1
0
13 Logic Switch~
5 839 906 0 1 11
0 10
0
0 0 21360 90
2 0V
-3 27 11 35
2 B0
-4 14 10 22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8862 0 0
2
44257.6 0
0
13 Logic Switch~
5 745 903 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-5 25 9 33
2 B3
-5 14 9 22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3202 0 0
2
44257.6 1
0
13 Logic Switch~
5 778 904 0 1 11
0 7
0
0 0 21360 90
2 0V
-5 26 9 34
2 B2
-5 14 9 22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5657 0 0
2
44257.6 0
0
13 Logic Switch~
5 481 895 0 1 11
0 12
0
0 0 21360 90
2 0V
-7 35 7 43
2 A1
-6 18 8 26
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3554 0 0
2
44257.6 1
0
13 Logic Switch~
5 515 897 0 1 11
0 11
0
0 0 21360 90
2 0V
-9 33 5 41
2 A0
-8 17 6 25
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4316 0 0
2
44257.6 0
0
13 Logic Switch~
5 447 897 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-7 32 7 40
2 A2
-6 18 8 26
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3739 0 0
2
44257.6 1
0
13 Logic Switch~
5 414 897 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-6 33 8 41
2 A3
-5 18 9 26
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7606 0 0
2
44257.6 0
0
13 Logic Switch~
5 415 630 0 10 11
0 32 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-5 -25 9 -17
2 S1
-31 -10 -17 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3741 0 0
2
44257.6 1
0
13 Logic Switch~
5 451 628 0 10 11
0 33 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 S0
14 -5 28 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
369 0 0
2
44257.6 0
0
13 Logic Switch~
5 198 306 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 C12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8773 0 0
2
44257.6 0
0
13 Logic Switch~
5 87 452 0 10 11
0 38 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-32 -5 -18 3
2 I0
19 4 33 12
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7981 0 0
2
44257.6 11
0
13 Logic Switch~
5 89 427 0 10 11
0 39 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-32 -5 -18 3
2 I1
18 3 32 11
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4205 0 0
2
44257.6 10
0
13 Logic Switch~
5 89 405 0 1 11
0 40
0
0 0 21360 0
2 0V
-32 -5 -18 3
2 I2
16 4 30 12
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3375 0 0
2
44257.6 9
0
13 Logic Switch~
5 88 385 0 10 11
0 45 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-32 -5 -18 3
2 I3
12 3 26 11
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
719 0 0
2
44257.6 8
0
13 Logic Switch~
5 89 364 0 1 11
0 44
0
0 0 21360 0
2 0V
-32 -5 -18 3
2 I4
15 -11 29 -3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3749 0 0
2
44257.6 7
0
13 Logic Switch~
5 91 340 0 10 11
0 43 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-32 -5 -18 3
2 I5
18 -10 32 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3871 0 0
2
44257.6 6
0
13 Logic Switch~
5 92 318 0 1 11
0 42
0
0 0 21360 0
2 0V
-32 -5 -18 3
2 I6
19 -12 33 -4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4393 0 0
2
44257.6 5
0
13 Logic Switch~
5 93 294 0 1 11
0 41
0
0 0 21360 0
2 0V
-32 -5 -18 3
2 I7
18 -12 32 -4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6229 0 0
2
44257.6 4
0
13 Logic Switch~
5 316 299 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 S2
-7 -31 7 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3757 0 0
2
44257.6 2
0
13 Logic Switch~
5 350 296 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 S1
-7 -31 7 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
352 0 0
2
44257.6 1
0
13 Logic Switch~
5 381 299 0 10 11
0 36 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 S0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3372 0 0
2
44257.6 0
0
13 Logic Switch~
5 587 193 0 10 11
0 46 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-32 -5 -18 3
1 C
24 -12 31 -4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4911 0 0
2
44257.6 0
0
13 Logic Switch~
5 586 101 0 1 11
0 47
0
0 0 21360 0
2 0V
-32 0 -18 8
1 S
26 -10 33 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7574 0 0
2
44257.6 0
0
13 Logic Switch~
5 113 174 0 1 11
0 50
0
0 0 21360 0
2 0V
-30 -7 -16 1
1 C
21 -11 28 -3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6601 0 0
2
44257.6 0
0
13 Logic Switch~
5 111 96 0 1 11
0 51
0
0 0 21360 0
2 0V
-33 -2 -19 6
1 S
23 -14 30 -6
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8531 0 0
2
44257.6 0
0
14 Logic Display~
6 596 521 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6532 0 0
2
44257.7 0
0
14 Logic Display~
6 632 518 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3621 0 0
2
44257.7 0
0
14 Logic Display~
6 662 520 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5174 0 0
2
44257.7 0
0
14 Logic Display~
6 697 517 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5452 0 0
2
44257.7 0
0
9 2-In XOR~
219 809 775 0 3 22
0 11 10 19
0
0 0 624 90
5 74F86
-18 -24 17 -16
3 U9D
-595 -255 -574 -247
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
3626 0 0
2
44257.6 0
0
9 2-In XOR~
219 677 774 0 3 22
0 12 9 23
0
0 0 624 90
5 74F86
-18 -24 17 -16
3 U9C
77 -496 98 -488
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
3806 0 0
2
44257.6 0
0
9 2-In XOR~
219 505 779 0 3 22
0 13 7 28
0
0 0 624 90
5 74F86
-18 -24 17 -16
3 U9B
255 -503 276 -495
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3389 0 0
2
44257.6 0
0
9 2-In XOR~
219 331 784 0 3 22
0 14 8 24
0
0 0 624 90
5 74F86
-18 -24 17 -16
3 U9A
415 -519 436 -511
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
9156 0 0
2
44257.6 0
0
9 Inverter~
13 912 773 0 2 22
0 11 22
0
0 0 624 90
5 74F04
-18 -19 17 -11
3 U8D
-700 -165 -679 -157
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 5 0
1 U
5810 0 0
2
44257.6 0
0
9 Inverter~
13 779 774 0 2 22
0 12 18
0
0 0 624 90
5 74F04
-18 -19 17 -11
3 U8C
-565 -185 -544 -177
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 5 0
1 U
8260 0 0
2
44257.6 0
0
9 Inverter~
13 615 778 0 2 22
0 13 31
0
0 0 624 90
5 74F04
-18 -19 17 -11
3 U8B
145 -523 166 -515
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 5 0
1 U
7286 0 0
2
44257.6 0
0
9 Inverter~
13 441 781 0 2 22
0 14 27
0
0 0 624 90
5 74F04
-18 -19 17 -11
3 U8A
-231 -251 -210 -243
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
3689 0 0
2
44257.6 0
0
8 2-In OR~
219 846 776 0 3 22
0 11 10 20
0
0 0 624 90
5 74F32
-18 -24 17 -16
3 U7D
-633 -206 -612 -198
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
4485 0 0
2
44257.6 0
0
8 2-In OR~
219 541 779 0 3 22
0 13 7 29
0
0 0 624 90
5 74F32
-18 -24 17 -16
3 U7C
219 -445 240 -437
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
4370 0 0
2
44257.6 0
0
8 2-In OR~
219 713 775 0 3 22
0 12 9 16
0
0 0 624 90
5 74F32
-18 -24 17 -16
3 U7B
-503 -233 -482 -225
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
7483 0 0
2
44257.6 0
0
8 2-In OR~
219 369 785 0 3 22
0 14 8 25
0
0 0 624 90
5 74F32
-18 -24 17 -16
3 U7A
-221 -267 -200 -259
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
4214 0 0
2
44257.6 0
0
9 2-In AND~
219 886 771 0 3 22
0 11 10 21
0
0 0 624 90
5 74F08
-18 -24 17 -16
3 U6D
-685 -192 -664 -184
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
9254 0 0
2
44257.6 0
0
9 2-In AND~
219 752 772 0 3 22
0 12 9 17
0
0 0 624 90
5 74F08
-18 -24 17 -16
3 U6C
4 -475 25 -467
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
7515 0 0
2
44257.6 0
0
9 2-In AND~
219 582 776 0 3 22
0 13 7 30
0
0 0 624 90
5 74F08
-18 -24 17 -16
3 U6B
-372 -223 -351 -215
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9241 0 0
2
44257.6 0
0
9 2-In AND~
219 411 781 0 3 22
0 14 8 26
0
0 0 624 90
5 74F08
-18 -24 17 -16
3 U6A
340 -496 361 -488
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3783 0 0
2
44257.6 0
0
7 74LS153
119 715 610 0 14 29
0 23 16 17 18 32 33 19 20 21
22 2 2 5 6
0
0 0 4848 90
6 74F153
-21 -60 21 -52
2 U5
-639 -22 -625 -14
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 0 0 0 0 0
1 U
5226 0 0
2
44257.6 0
0
7 74LS153
119 572 612 0 14 29
0 24 25 26 27 32 33 28 29 30
31 2 2 3 4
0
0 0 4848 90
6 74F153
-21 -60 21 -52
2 U4
-495 -49 -481 -41
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 0 0 0 0 0
1 U
6496 0 0
2
44257.6 0
0
7 74LS151
20 251 370 0 14 29
0 41 42 43 44 45 40 39 38 15
34 35 36 37 15
0
0 0 4848 0
6 74F151
-21 -60 21 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 0 0 0 0
1 U
6819 0 0
2
44257.6 12
0
14 Logic Display~
6 341 389 0 1 2
10 37
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L5
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6832 0 0
2
44257.6 3
0
14 Logic Display~
6 814 168 0 1 2
10 53
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7222 0 0
2
44257.6 0
0
14 Logic Display~
6 813 94 0 1 2
10 52
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4676 0 0
2
44257.6 0
0
14 Logic Display~
6 372 146 0 1 2
10 49
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9334 0 0
2
44257.6 0
0
14 Logic Display~
6 372 88 0 1 2
10 48
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4758 0 0
2
44257.6 0
0
10 2-In NAND~
219 247 105 0 3 22
0 51 49 48
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
6695 0 0
2
5.89975e-315 5.32571e-315
0
10 2-In NAND~
219 247 165 0 3 22
0 48 50 49
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
8212 0 0
2
5.89975e-315 5.30499e-315
0
9 2-In NOR~
219 702 111 0 3 22
0 47 53 52
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U1B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3922 0 0
2
5.89975e-315 5.26354e-315
0
9 2-In NOR~
219 704 185 0 3 22
0 52 46 53
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
7610 0 0
2
5.89975e-315 0
0
82
11 0 2 0 0 4096 0 49 0 0 4 3
537 579
537 570
538 570
12 0 2 0 0 0 0 49 0 0 4 3
618 579
618 570
619 570
11 0 2 0 0 0 0 48 0 0 4 3
680 577
680 570
679 570
1 12 2 0 0 4224 0 1 48 0 0 3
510 570
761 570
761 577
1 13 3 0 0 8336 0 28 49 0 0 4
596 539
596 544
555 544
555 585
1 14 4 0 0 8320 0 29 49 0 0 4
632 536
632 560
600 560
600 585
1 13 5 0 0 8320 0 30 48 0 0 4
662 538
662 559
698 559
698 583
1 14 6 0 0 8320 0 31 48 0 0 4
697 535
697 544
743 544
743 583
2 0 7 0 0 4096 0 46 0 0 19 2
590 797
590 853
2 0 7 0 0 4096 0 41 0 0 19 2
553 795
553 853
2 0 8 0 0 4096 0 47 0 0 20 2
419 802
419 859
2 0 8 0 0 4096 0 43 0 0 20 2
381 801
381 859
2 0 9 0 0 4096 0 42 0 0 14 2
725 791
725 847
0 2 9 0 0 4096 0 0 45 18 0 3
689 847
760 847
760 793
2 0 10 0 0 4096 0 40 0 0 16 2
858 792
858 845
0 2 10 0 0 4096 0 0 44 17 0 3
821 845
894 845
894 792
2 1 10 0 0 4224 0 32 3 0 0 4
821 794
821 886
840 886
840 893
2 1 9 0 0 8320 0 33 2 0 0 4
689 793
689 884
811 884
811 891
2 1 7 0 0 8320 0 34 5 0 0 4
517 798
517 853
779 853
779 891
2 1 8 0 0 8320 0 35 4 0 0 4
343 803
343 859
746 859
746 890
1 0 11 0 0 4096 0 40 0 0 23 2
840 792
840 823
1 0 11 0 0 0 0 44 0 0 23 2
876 792
876 823
0 1 11 0 0 4096 0 0 36 24 0 3
803 823
915 823
915 791
1 1 11 0 0 8320 0 7 32 0 0 4
516 884
516 873
803 873
803 794
1 0 12 0 0 4096 0 45 0 0 27 2
742 793
742 824
1 0 12 0 0 4096 0 42 0 0 27 2
707 791
707 824
0 1 12 0 0 4096 0 0 37 28 0 3
671 824
782 824
782 792
1 1 12 0 0 8320 0 33 6 0 0 4
671 793
671 867
482 867
482 882
1 0 13 0 0 4096 0 46 0 0 31 2
572 797
572 833
1 0 13 0 0 4096 0 41 0 0 31 2
535 795
535 833
0 1 13 0 0 4224 0 0 38 32 0 3
499 833
618 833
618 796
1 1 13 0 0 0 0 34 8 0 0 4
499 798
499 834
448 834
448 884
1 0 14 0 0 4096 0 47 0 0 35 2
401 802
401 833
1 0 14 0 0 0 0 43 0 0 35 4
363 801
363 828
364 828
364 833
0 1 14 0 0 4224 0 0 39 36 0 3
325 833
444 833
444 799
1 1 14 0 0 0 0 9 35 0 0 4
415 884
415 871
325 871
325 803
9 1 15 0 0 12416 0 50 12 0 0 4
289 343
293 343
293 306
210 306
2 3 16 0 0 4224 0 48 42 0 0 4
689 647
689 744
716 744
716 745
3 3 17 0 0 4224 0 48 45 0 0 4
698 647
698 735
751 735
751 748
4 2 18 0 0 4224 0 48 37 0 0 4
707 647
707 729
782 729
782 756
7 3 19 0 0 8320 0 48 32 0 0 4
734 647
734 720
812 720
812 745
8 3 20 0 0 8320 0 48 40 0 0 4
743 647
743 709
849 709
849 746
9 3 21 0 0 8320 0 48 44 0 0 4
752 647
752 697
885 697
885 747
10 2 22 0 0 8320 0 48 36 0 0 4
761 647
761 686
915 686
915 755
1 3 23 0 0 4224 0 48 33 0 0 2
680 647
680 744
1 3 24 0 0 8320 0 49 35 0 0 4
537 649
537 690
334 690
334 754
2 3 25 0 0 8320 0 49 43 0 0 4
546 649
546 702
372 702
372 755
3 3 26 0 0 8320 0 49 47 0 0 4
555 649
555 711
410 711
410 757
4 2 27 0 0 8320 0 49 39 0 0 4
564 649
564 720
444 720
444 763
7 3 28 0 0 8320 0 49 34 0 0 4
591 649
591 731
508 731
508 749
8 3 29 0 0 4224 0 49 41 0 0 4
600 649
600 738
544 738
544 749
9 3 30 0 0 4224 0 49 46 0 0 4
609 649
609 746
581 746
581 752
10 2 31 0 0 4224 0 49 38 0 0 2
618 649
618 760
0 1 32 0 0 8320 0 0 10 56 0 4
658 660
658 681
415 681
415 642
0 1 33 0 0 8320 0 0 11 57 0 4
645 655
645 672
451 672
451 640
5 5 32 0 0 0 0 49 48 0 0 4
573 649
573 660
716 660
716 647
6 6 33 0 0 0 0 49 48 0 0 4
582 649
582 655
725 655
725 647
9 14 15 0 0 128 0 50 50 0 0 4
289 343
302 343
302 406
289 406
10 1 34 0 0 8320 0 50 21 0 0 3
283 352
316 352
316 311
11 1 35 0 0 4224 0 50 22 0 0 3
283 361
350 361
350 308
12 1 36 0 0 4224 0 50 23 0 0 3
283 370
381 370
381 311
13 1 37 0 0 4224 0 50 51 0 0 4
283 397
318 397
318 393
325 393
8 1 38 0 0 4224 0 50 13 0 0 4
219 406
139 406
139 452
99 452
7 1 39 0 0 4224 0 50 14 0 0 4
219 397
129 397
129 427
101 427
6 1 40 0 0 4224 0 50 15 0 0 4
219 388
119 388
119 405
101 405
1 1 41 0 0 4224 0 50 20 0 0 4
219 343
137 343
137 294
105 294
2 1 42 0 0 4224 0 50 19 0 0 4
219 352
128 352
128 318
104 318
3 1 43 0 0 4224 0 50 18 0 0 4
219 361
122 361
122 340
103 340
4 1 44 0 0 4224 0 50 17 0 0 4
219 370
110 370
110 364
101 364
5 1 45 0 0 4224 0 50 16 0 0 4
219 379
110 379
110 385
100 385
1 2 46 0 0 8320 0 24 59 0 0 3
599 193
599 194
691 194
1 1 47 0 0 8320 0 25 58 0 0 3
598 101
598 102
689 102
0 1 48 0 0 8320 0 0 57 76 0 5
305 105
305 128
159 128
159 156
223 156
2 0 49 0 0 12416 0 56 0 0 75 5
223 114
174 114
174 138
305 138
305 165
3 1 49 0 0 0 0 57 54 0 0 3
274 165
372 165
372 164
3 1 48 0 0 0 0 56 55 0 0 4
274 105
305 105
305 106
372 106
1 2 50 0 0 4224 0 26 57 0 0 2
125 174
223 174
1 1 51 0 0 4224 0 27 56 0 0 2
123 96
223 96
1 0 52 0 0 12416 0 59 0 0 82 5
691 176
646 176
646 141
764 141
764 111
2 0 53 0 0 12416 0 58 0 0 81 5
689 120
627 120
627 155
767 155
767 185
3 1 53 0 0 0 0 59 52 0 0 3
743 185
814 185
814 186
3 1 52 0 0 0 0 58 53 0 0 3
741 111
813 111
813 112
66
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
777 830 812 851
786 836 802 851
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
794 786 829 807
803 793 819 808
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
805 722 840 743
814 729 830 744
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
671 794 694 815
678 801 686 816
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
643 822 676 843
651 829 667 844
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
655 728 680 749
663 735 671 750
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
488 734 513 755
496 741 504 756
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
499 797 526 818
508 804 516 819
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
474 787 501 808
483 794 491 809
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
330 732 357 753
339 739 347 754
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
338 801 363 822
346 807 354 822
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
304 809 331 830
313 815 321 830
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
845 722 880 743
854 729 870 744
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
832 786 867 807
841 793 857 808
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
825 818 860 839
834 824 850 839
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
712 730 737 751
720 737 728 752
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
709 788 732 809
716 795 724 810
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
691 820 724 841
699 827 715 842
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
544 734 569 755
552 741 560 756
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
523 828 550 849
532 835 540 850
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
534 790 561 811
543 797 551 812
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
366 733 393 754
375 740 383 755
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
377 796 402 817
385 802 393 817
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
350 828 377 849
359 834 367 849
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
879 723 914 744
888 730 904 745
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
862 820 897 841
871 826 887 841
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
868 786 903 807
877 793 893 808
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
747 728 772 749
755 735 763 750
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
726 820 759 841
734 827 750 842
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
744 787 767 808
751 794 759 809
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
584 741 609 762
592 748 600 763
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
559 828 586 849
568 835 576 850
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
572 792 599 813
581 799 589 814
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
406 732 433 753
415 739 423 754
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
388 827 415 848
397 833 405 848
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
414 796 439 817
422 802 430 817
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
911 724 936 745
919 731 927 746
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
911 803 938 824
920 809 928 824
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
776 738 803 759
785 745 793 760
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
776 795 801 816
784 802 792 817
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
613 737 640 758
622 743 630 758
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
613 796 640 817
622 803 630 818
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
439 736 464 757
447 742 455 757
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
442 789 467 810
450 796 458 811
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
822 640 885 664
829 645 877 661
6 3-X-OR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
821 616 868 640
828 622 860 638
4 2-OR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
821 596 876 620
828 602 868 618
5 1-AND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
822 574 877 598
829 579 869 595
5 0-NOT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
665 192 690 213
673 199 681 214
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
663 155 690 176
672 162 680 177
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
763 186 790 207
772 193 780 208
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
664 115 691 136
673 121 681 136
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
663 75 690 96
672 82 680 97
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
768 87 795 108
777 93 785 108
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
321 146 346 167
329 153 337 168
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
186 168 211 189
194 175 202 190
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
185 134 210 155
193 141 201 156
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
317 79 344 100
326 86 334 101
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
186 93 211 114
194 99 202 114
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
186 72 213 93
195 78 203 93
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
828 75 865 99
838 83 854 99
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
381 124 418 148
391 132 407 148
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
838 162 867 186
848 170 856 186
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
832 89 861 113
842 97 850 113
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
385 140 414 164
395 148 403 164
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
381 80 410 104
391 88 399 104
1 Q
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
