CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
190 330 30 110 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
75
13 Logic Switch~
5 1049 848 0 1 11
0 3
0
0 0 21360 90
2 0V
-4 27 10 35
2 B1
-5 16 9 24
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5179 0 0
2
44279.9 0
0
13 Logic Switch~
5 1080 849 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-3 27 11 35
2 B0
-4 14 10 22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3593 0 0
2
44279.9 1
0
13 Logic Switch~
5 983 850 0 1 11
0 5
0
0 0 21360 90
2 0V
-5 25 9 33
2 B3
-5 14 9 22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3928 0 0
2
44279.9 2
0
13 Logic Switch~
5 1019 849 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-5 26 9 34
2 B2
-5 14 9 22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
363 0 0
2
44279.9 3
0
13 Logic Switch~
5 770 852 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-6 33 8 41
2 A3
-5 18 9 26
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8132 0 0
2
44279.9 4
0
13 Logic Switch~
5 801 850 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-7 32 7 40
2 A2
-6 18 8 26
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
65 0 0
2
44279.9 5
0
13 Logic Switch~
5 867 849 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-9 33 5 41
2 A0
-8 17 6 25
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6609 0 0
2
44279.9 6
0
13 Logic Switch~
5 836 849 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
-7 35 7 43
2 A1
-6 18 8 26
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8995 0 0
2
44279.9 7
0
13 Logic Switch~
5 738 551 0 1 11
0 26
0
0 0 21360 0
2 0V
-31 -4 -17 4
3 C15
872 -292 893 -284
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3918 0 0
2
44279.9 8
0
13 Logic Switch~
5 820 405 0 1 11
0 39
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 Cin
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7519 0 0
2
5.89977e-315 0
0
13 Logic Switch~
5 791 405 0 10 11
0 33 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 S0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
377 0 0
2
5.89977e-315 5.26354e-315
0
13 Logic Switch~
5 765 405 0 1 11
0 32
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 S1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8816 0 0
2
5.89977e-315 5.30499e-315
0
13 Logic Switch~
5 731 405 0 10 11
0 38 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 S
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3877 0 0
2
5.89977e-315 5.32571e-315
0
9 Inverter~
13 828 747 0 2 22
0 8 14
0
0 0 624 90
5 74F04
-18 -19 17 -11
3 U4E
712 -491 733 -483
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 4 0
1 U
926 0 0
2
5.89977e-315 0
0
9 Inverter~
13 692 747 0 2 22
0 9 10
0
0 0 624 90
5 74F04
-18 -19 17 -11
4 U12C
853 -491 881 -483
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 11 0
1 U
7262 0 0
2
5.89977e-315 0
0
9 2-In XOR~
219 933 746 0 3 22
0 8 4 17
0
0 0 624 90
5 74F86
-18 -24 17 -16
4 U13D
939 -568 967 -560
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 12 0
1 U
5267 0 0
2
5.89977e-315 5.26354e-315
0
9 2-In XOR~
219 770 1199 0 3 22
0 75 76 77
0
0 0 624 90
5 74F86
-18 -24 17 -16
4 U13C
939 -568 967 -560
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 12 0
1 U
8838 0 0
2
5.89977e-315 0
0
9 2-In XOR~
219 652 1139 0 3 22
0 78 79 80
0
0 0 624 90
5 74F86
-18 -24 17 -16
4 U13B
939 -568 967 -560
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 12 0
1 U
7159 0 0
2
5.89977e-315 0
0
9 2-In XOR~
219 794 745 0 3 22
0 9 5 13
0
0 0 624 90
5 74F86
-18 -24 17 -16
4 U13A
939 -568 967 -560
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
5812 0 0
2
5.89977e-315 0
0
8 2-In OR~
219 1041 747 0 3 22
0 7 3 19
0
0 0 624 90
5 74F32
-18 -24 17 -16
4 U20A
845 -443 873 -435
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 17 0
1 U
331 0 0
2
5.89977e-315 5.26354e-315
0
8 2-In OR~
219 1180 745 0 3 22
0 6 2 24
0
0 0 624 90
5 74F32
-18 -24 17 -16
4 U17D
845 -443 873 -435
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
9604 0 0
2
5.89977e-315 0
0
8 2-In OR~
219 896 749 0 3 22
0 8 4 16
0
0 0 624 90
5 74F32
-18 -24 17 -16
4 U17B
845 -443 873 -435
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
7518 0 0
2
5.89977e-315 0
0
9 2-In AND~
219 862 744 0 3 22
0 8 4 15
0
0 0 624 90
5 74F08
-18 -24 17 -16
4 U19A
850 -563 878 -555
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
4832 0 0
2
5.89977e-315 5.26354e-315
0
9 2-In AND~
219 1148 742 0 3 22
0 6 2 23
0
0 0 624 90
5 74F08
-18 -24 17 -16
4 U18C
850 -563 878 -555
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
6798 0 0
2
5.89977e-315 0
0
9 2-In AND~
219 1008 745 0 3 22
0 7 3 20
0
0 0 624 90
5 74F08
-18 -24 17 -16
4 U18B
850 -563 878 -555
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
3336 0 0
2
5.89977e-315 0
0
9 2-In AND~
219 726 744 0 3 22
0 9 5 11
0
0 0 624 90
5 74F08
-18 -24 17 -16
4 U18A
850 -563 878 -555
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
8370 0 0
2
5.89977e-315 0
0
8 2-In OR~
219 757 747 0 3 22
0 9 5 12
0
0 0 624 90
5 74F32
-18 -24 17 -16
4 U17A
845 -443 873 -435
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
3910 0 0
2
5.89977e-315 0
0
14 Logic Display~
6 961 419 0 1 2
10 27
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
316 0 0
2
44279.9 9
0
14 Logic Display~
6 1015 422 0 1 2
10 28
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
536 0 0
2
44279.9 10
0
14 Logic Display~
6 1035 422 0 1 2
10 29
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4460 0 0
2
44279.9 11
0
14 Logic Display~
6 1059 422 0 1 2
10 30
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3260 0 0
2
44279.9 12
0
14 Logic Display~
6 1081 422 0 1 2
10 31
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5156 0 0
2
44279.9 13
0
7 74LS153
119 898 589 0 14 29
0 10 11 12 13 32 33 14 15 16
17 26 26 34 35
0
0 0 4848 90
6 74F153
-21 -60 21 -52
3 U16
692 -272 713 -264
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 0 1 0 0 0
1 U
3133 0 0
2
44279.9 14
0
7 74LS153
119 1018 590 0 14 29
0 21 20 19 18 32 33 22 23 24
25 26 26 36 37
0
0 0 4848 90
6 74F153
-21 -60 21 -52
3 U15
518 -270 539 -262
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 0 1 0 0 0
1 U
5523 0 0
2
44279.9 15
0
9 Inverter~
13 974 748 0 2 22
0 7 21
0
0 0 624 90
5 74F04
-18 -19 17 -11
3 U4F
572 -497 593 -489
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 4 0
1 U
3746 0 0
2
44279.9 16
0
9 Inverter~
13 1113 745 0 2 22
0 6 22
0
0 0 624 90
5 74F04
-18 -19 17 -11
3 U4E
419 -486 440 -478
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 4 0
1 U
5668 0 0
2
44279.9 17
0
9 2-In XOR~
219 1078 744 0 3 22
0 7 3 18
0
0 0 624 90
5 74F86
-18 -24 17 -16
4 U11B
612 -557 640 -549
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
5368 0 0
2
44279.9 18
0
9 2-In XOR~
219 1216 742 0 3 22
0 6 2 25
0
0 0 624 90
5 74F86
-18 -24 17 -16
4 U11A
418 -434 446 -426
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
8293 0 0
2
44279.9 19
0
7 74LS257
147 881 475 0 14 29
0 38 34 40 35 41 36 42 37 43
26 28 29 30 31
0
0 0 4848 0
6 74F257
-21 -60 21 -52
3 U10
726 -155 747 -147
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3232 0 0
2
44279.9 20
0
9 Inverter~
13 285 724 0 2 22
0 5 51
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4D
1355 -408 1376 -400
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 4 0
1 U
6644 0 0
2
44279.9 21
0
8 2-In OR~
219 414 713 0 3 22
0 53 52 48
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U8D
1177 -393 1198 -385
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
4978 0 0
2
44279.9 22
0
9 2-In AND~
219 356 732 0 3 22
0 51 32 52
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U9D
1273 -432 1294 -424
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
9207 0 0
2
44279.9 23
0
9 2-In AND~
219 361 696 0 3 22
0 5 33 53
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U9C
1272 -358 1293 -350
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
6998 0 0
2
44279.9 24
0
8 2-In OR~
219 629 743 0 3 22
0 49 50 27
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U8C
965 -423 986 -415
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
3175 0 0
2
44279.9 25
0
9 2-In AND~
219 579 725 0 3 22
0 47 44 49
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U9B
1022 -403 1043 -395
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
3378 0 0
2
44279.9 26
0
9 2-In AND~
219 506 752 0 3 22
0 48 9 50
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U9A
1061 -431 1082 -423
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
922 0 0
2
44279.9 27
0
9 2-In XOR~
219 632 693 0 3 22
0 44 47 40
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6D
966 -368 987 -360
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
6891 0 0
2
44279.9 28
0
9 2-In XOR~
219 500 703 0 3 22
0 9 48 47
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6C
1077 -372 1098 -364
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
5407 0 0
2
44279.9 29
0
9 Inverter~
13 286 624 0 2 22
0 4 58
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4C
1355 -408 1376 -400
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
7349 0 0
2
44279.9 30
0
8 2-In OR~
219 415 613 0 3 22
0 60 59 55
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U8B
1177 -393 1198 -385
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
3919 0 0
2
44279.9 31
0
9 2-In AND~
219 357 632 0 3 22
0 58 32 59
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7D
1273 -432 1294 -424
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
9747 0 0
2
44279.9 32
0
9 2-In AND~
219 362 596 0 3 22
0 4 33 60
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7C
1272 -358 1293 -350
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
5310 0 0
2
44279.9 33
0
8 2-In OR~
219 630 643 0 3 22
0 56 57 44
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U8A
1027 -407 1048 -399
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
4318 0 0
2
44279.9 34
0
9 2-In AND~
219 580 625 0 3 22
0 54 45 56
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7B
963 -385 984 -377
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
3917 0 0
2
44279.9 35
0
9 2-In AND~
219 507 652 0 3 22
0 55 8 57
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7A
1061 -431 1082 -423
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
7930 0 0
2
44279.9 36
0
9 2-In XOR~
219 633 593 0 3 22
0 45 54 41
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6B
932 -333 953 -325
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
6128 0 0
2
44279.9 37
0
9 2-In XOR~
219 501 603 0 3 22
0 8 55 54
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6A
1077 -372 1098 -364
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
7346 0 0
2
44279.9 38
0
9 Inverter~
13 285 525 0 2 22
0 3 65
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4B
1355 -408 1376 -400
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
8577 0 0
2
44279.9 39
0
8 2-In OR~
219 414 514 0 3 22
0 67 66 62
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3D
1177 -393 1198 -385
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3372 0 0
2
44279.9 40
0
9 2-In AND~
219 356 533 0 3 22
0 65 32 66
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5D
1273 -432 1294 -424
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3741 0 0
2
44279.9 41
0
9 2-In AND~
219 361 497 0 3 22
0 3 33 67
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5C
1272 -358 1293 -350
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
5813 0 0
2
44279.9 42
0
8 2-In OR~
219 629 544 0 3 22
0 63 64 45
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3C
1029 -398 1050 -390
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3213 0 0
2
44279.9 43
0
9 2-In AND~
219 579 526 0 3 22
0 61 46 63
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5B
963 -385 984 -377
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3694 0 0
2
44279.9 44
0
9 2-In AND~
219 506 553 0 3 22
0 62 7 64
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5A
1061 -431 1082 -423
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
4327 0 0
2
44279.9 45
0
9 2-In XOR~
219 632 494 0 3 22
0 46 61 42
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1D
932 -333 953 -325
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
8800 0 0
2
44279.9 46
0
9 2-In XOR~
219 500 504 0 3 22
0 7 62 61
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1C
1077 -372 1098 -364
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3406 0 0
2
44279.9 47
0
9 2-In XOR~
219 499 402 0 3 22
0 6 69 68
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1A
1077 -372 1098 -364
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
6455 0 0
2
44279.9 48
0
9 2-In XOR~
219 631 392 0 3 22
0 39 68 43
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1B
932 -333 953 -325
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9319 0 0
2
44279.9 49
0
9 2-In AND~
219 505 451 0 3 22
0 69 6 71
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2A
1061 -431 1082 -423
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3172 0 0
2
44279.9 50
0
9 2-In AND~
219 578 424 0 3 22
0 68 39 70
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2B
963 -385 984 -377
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
38 0 0
2
44279.9 51
0
8 2-In OR~
219 628 442 0 3 22
0 70 71 46
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3A
872 -400 893 -392
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
376 0 0
2
44279.9 52
0
9 2-In AND~
219 360 395 0 3 22
0 2 33 74
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2C
1272 -358 1293 -350
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
6666 0 0
2
44279.9 53
0
9 2-In AND~
219 355 431 0 3 22
0 72 32 73
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2D
1273 -432 1294 -424
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
9365 0 0
2
44279.9 54
0
8 2-In OR~
219 413 412 0 3 22
0 74 73 69
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3B
1177 -393 1198 -385
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3251 0 0
2
44279.9 55
0
9 Inverter~
13 284 423 0 2 22
0 2 72
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4A
1355 -408 1376 -400
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
5481 0 0
2
44279.9 56
0
135
0 0 2 0 0 4224 0 0 0 9 129 4
1081 828
208 828
208 386
262 386
0 0 3 0 0 12416 0 0 0 118 10 4
263 488
247 488
247 824
1030 824
0 0 4 0 0 12416 0 0 0 107 11 4
264 587
241 587
241 819
1000 819
0 0 5 0 0 12416 0 0 0 96 12 4
263 687
219 687
219 815
734 815
0 0 6 0 0 4224 0 0 0 13 62 4
871 810
224 810
224 460
454 460
0 0 7 0 0 4224 0 0 0 14 61 4
837 805
229 805
229 562
451 562
0 0 8 0 0 4224 0 0 0 15 60 4
812 800
233 800
233 661
452 661
0 0 9 0 0 8320 0 0 0 59 16 3
453 761
453 774
695 774
0 1 2 0 0 0 0 0 2 21 0 5
1156 787
1126 787
1126 809
1081 809
1081 836
1 0 3 0 0 0 0 1 0 0 22 6
1050 835
1050 834
1030 834
1030 809
1016 809
1016 788
0 1 4 0 0 0 0 0 4 23 0 6
943 788
943 809
1000 809
1000 833
1020 833
1020 836
0 1 5 0 0 0 0 0 3 24 0 4
734 785
734 833
984 833
984 837
1 0 6 0 0 0 0 7 0 0 49 7
868 836
868 810
871 810
871 804
1115 804
1115 774
1116 774
0 1 7 0 0 0 0 0 8 50 0 4
977 776
977 800
837 800
837 836
1 0 8 0 0 0 0 6 0 0 51 4
802 837
812 837
812 776
831 776
1 0 9 0 0 0 0 5 0 0 52 4
771 839
771 838
695 838
695 774
2 0 2 0 0 0 0 21 0 0 21 2
1192 761
1192 787
2 0 3 0 0 0 0 20 0 0 22 2
1053 763
1053 788
2 0 4 0 0 0 0 22 0 0 23 2
908 765
908 788
2 0 5 0 0 0 0 27 0 0 24 2
769 763
769 787
2 2 2 0 0 0 0 24 38 0 0 4
1156 763
1156 787
1228 787
1228 761
2 2 3 0 0 0 0 25 37 0 0 4
1016 766
1016 788
1090 788
1090 763
2 2 4 0 0 0 0 23 16 0 0 4
870 765
870 788
945 788
945 765
2 2 5 0 0 0 0 26 19 0 0 4
734 765
734 787
806 787
806 764
2 1 10 0 0 8320 0 15 33 0 0 4
695 729
695 667
863 667
863 626
3 2 11 0 0 8320 0 26 33 0 0 4
725 720
725 673
872 673
872 626
3 3 12 0 0 8320 0 27 33 0 0 4
760 717
760 677
881 677
881 626
3 4 13 0 0 8320 0 19 33 0 0 4
797 715
797 683
890 683
890 626
2 7 14 0 0 8320 0 14 33 0 0 4
831 729
831 690
917 690
917 626
3 8 15 0 0 12416 0 23 33 0 0 4
861 720
861 696
926 696
926 626
3 9 16 0 0 12416 0 22 33 0 0 4
899 719
899 702
935 702
935 626
3 10 17 0 0 12416 0 16 33 0 0 4
936 716
936 708
944 708
944 626
3 4 18 0 0 8320 0 37 34 0 0 4
1081 714
1081 685
1010 685
1010 627
3 3 19 0 0 12416 0 20 34 0 0 4
1044 717
1044 693
1001 693
1001 627
3 2 20 0 0 12416 0 25 34 0 0 4
1007 721
1007 699
992 699
992 627
2 1 21 0 0 12416 0 35 34 0 0 4
977 730
977 708
983 708
983 627
2 7 22 0 0 8320 0 36 34 0 0 4
1116 727
1116 675
1037 675
1037 627
3 8 23 0 0 8320 0 24 34 0 0 4
1147 718
1147 668
1046 668
1046 627
3 9 24 0 0 8320 0 21 34 0 0 4
1183 715
1183 658
1055 658
1055 627
3 10 25 0 0 8320 0 38 34 0 0 4
1219 712
1219 650
1064 650
1064 627
1 0 6 0 0 0 0 21 0 0 49 2
1174 761
1174 775
1 0 6 0 0 0 0 24 0 0 49 2
1138 763
1138 775
1 0 7 0 0 0 0 20 0 0 50 2
1035 763
1035 776
1 0 7 0 0 0 0 25 0 0 50 2
998 766
998 776
1 0 8 0 0 0 0 22 0 0 51 2
890 765
890 776
1 0 8 0 0 0 0 23 0 0 51 2
852 765
852 776
1 0 9 0 0 0 0 27 0 0 52 2
751 763
751 774
1 0 9 0 0 0 0 26 0 0 52 2
716 765
716 774
1 1 6 0 0 0 0 36 38 0 0 4
1116 763
1116 775
1210 775
1210 761
1 1 7 0 0 0 0 35 37 0 0 4
977 766
977 776
1072 776
1072 763
1 1 8 0 0 0 0 14 16 0 0 4
831 765
831 776
927 776
927 765
1 1 9 0 0 0 0 15 19 0 0 4
695 765
695 774
788 774
788 764
11 0 26 0 0 4096 0 33 0 0 72 3
863 556
863 550
862 550
1 3 27 0 0 8320 0 28 44 0 0 5
961 437
961 631
678 631
678 743
662 743
11 1 28 0 0 4224 0 39 29 0 0 3
913 457
1015 457
1015 440
12 1 29 0 0 4224 0 39 30 0 0 3
913 475
1035 475
1035 440
13 1 30 0 0 4224 0 39 31 0 0 3
913 493
1059 493
1059 440
14 1 31 0 0 4224 0 39 32 0 0 3
913 511
1081 511
1081 440
1 2 9 0 0 0 0 48 46 0 0 4
484 694
453 694
453 761
482 761
1 2 8 0 0 0 0 57 55 0 0 4
485 594
452 594
452 661
483 661
1 2 7 0 0 0 0 66 64 0 0 4
484 495
451 495
451 562
482 562
1 2 6 0 0 0 0 67 69 0 0 4
483 393
454 393
454 460
481 460
0 0 32 0 0 8320 0 0 0 85 73 4
237 741
237 792
966 792
966 655
11 0 26 0 0 4096 0 34 0 0 72 3
983 557
983 550
985 550
12 0 26 0 0 0 0 33 0 0 72 3
944 556
944 550
943 550
0 0 33 0 0 8336 0 0 0 88 74 4
214 705
214 796
959 796
959 645
13 2 34 0 0 12416 0 33 39 0 0 5
881 562
881 556
799 556
799 448
849 448
14 4 35 0 0 8320 0 33 39 0 0 5
926 562
926 544
807 544
807 466
849 466
13 6 36 0 0 8320 0 34 39 0 0 5
1001 563
1001 537
814 537
814 484
849 484
14 8 37 0 0 8320 0 34 39 0 0 5
1046 563
1046 532
820 532
820 502
849 502
10 0 26 0 0 8192 0 39 0 0 72 3
843 520
839 520
839 550
1 12 26 0 0 8320 0 9 34 0 0 4
750 551
750 550
1064 550
1064 557
0 1 32 0 0 0 0 0 12 75 0 4
978 640
978 655
765 655
765 417
0 1 33 0 0 0 0 0 11 76 0 4
959 635
959 645
791 645
791 417
5 5 32 0 0 0 0 33 34 0 0 4
899 626
899 640
1019 640
1019 627
6 6 33 0 0 0 0 33 34 0 0 4
908 626
908 635
1028 635
1028 627
1 1 38 0 0 8320 0 13 39 0 0 3
731 417
731 439
849 439
1 0 39 0 0 12416 0 10 0 0 125 5
820 417
907 417
907 366
537 366
537 383
3 3 40 0 0 8320 0 47 39 0 0 4
665 693
687 693
687 457
849 457
3 5 41 0 0 12416 0 56 39 0 0 4
666 593
675 593
675 475
849 475
3 7 42 0 0 12416 0 65 39 0 0 4
665 494
680 494
680 493
849 493
3 9 43 0 0 12416 0 68 39 0 0 4
664 392
681 392
681 511
849 511
2 0 32 0 0 0 0 51 0 0 85 2
333 641
237 641
2 0 32 0 0 0 0 60 0 0 85 2
332 542
237 542
2 2 32 0 0 0 0 73 42 0 0 4
331 440
237 440
237 741
332 741
2 0 33 0 0 0 0 52 0 0 88 2
338 605
214 605
2 0 33 0 0 0 0 61 0 0 88 2
337 506
214 506
2 2 33 0 0 0 0 72 43 0 0 4
336 404
214 404
214 705
337 705
3 0 44 0 0 12416 0 53 0 0 92 5
663 643
669 643
669 669
538 669
538 684
3 0 45 0 0 12416 0 62 0 0 103 5
662 544
670 544
670 568
539 568
539 584
3 0 46 0 0 12416 0 71 0 0 114 5
661 442
669 442
669 471
538 471
538 485
1 2 44 0 0 0 0 47 45 0 0 4
616 684
538 684
538 734
555 734
0 1 47 0 0 4096 0 0 45 99 0 3
548 703
548 716
555 716
3 0 48 0 0 4096 0 41 0 0 95 3
447 713
476 713
476 712
2 1 48 0 0 8320 0 48 46 0 0 4
484 712
476 712
476 743
482 743
1 1 5 0 0 0 0 43 40 0 0 4
337 687
263 687
263 724
270 724
3 1 49 0 0 12416 0 45 44 0 0 4
600 725
606 725
606 734
616 734
3 2 50 0 0 4224 0 46 44 0 0 2
527 752
616 752
3 2 47 0 0 4224 0 48 47 0 0 3
533 703
616 703
616 702
2 1 51 0 0 4224 0 40 42 0 0 4
306 724
329 724
329 723
332 723
3 2 52 0 0 12416 0 42 41 0 0 4
377 732
388 732
388 722
401 722
3 1 53 0 0 12416 0 43 41 0 0 4
382 696
389 696
389 704
401 704
1 2 45 0 0 0 0 56 54 0 0 4
617 584
539 584
539 634
556 634
0 1 54 0 0 4096 0 0 54 110 0 3
549 603
549 616
556 616
3 0 55 0 0 4096 0 50 0 0 106 3
448 613
477 613
477 612
2 1 55 0 0 8320 0 57 55 0 0 4
485 612
477 612
477 643
483 643
1 1 4 0 0 0 0 52 49 0 0 4
338 587
264 587
264 624
271 624
3 1 56 0 0 12416 0 54 53 0 0 4
601 625
607 625
607 634
617 634
3 2 57 0 0 4224 0 55 53 0 0 2
528 652
617 652
3 2 54 0 0 4224 0 57 56 0 0 3
534 603
617 603
617 602
2 1 58 0 0 4224 0 49 51 0 0 4
307 624
330 624
330 623
333 623
3 2 59 0 0 12416 0 51 50 0 0 4
378 632
389 632
389 622
402 622
3 1 60 0 0 12416 0 52 50 0 0 4
383 596
390 596
390 604
402 604
1 2 46 0 0 0 0 65 63 0 0 4
616 485
538 485
538 535
555 535
0 1 61 0 0 4096 0 0 63 121 0 3
548 504
548 517
555 517
3 0 62 0 0 4096 0 59 0 0 117 3
447 514
476 514
476 513
2 1 62 0 0 8320 0 66 64 0 0 4
484 513
476 513
476 544
482 544
1 1 3 0 0 0 0 61 58 0 0 4
337 488
263 488
263 525
270 525
3 1 63 0 0 12416 0 63 62 0 0 4
600 526
606 526
606 535
616 535
3 2 64 0 0 4224 0 64 62 0 0 2
527 553
616 553
3 2 61 0 0 4224 0 66 65 0 0 3
533 504
616 504
616 503
2 1 65 0 0 4224 0 58 60 0 0 4
306 525
329 525
329 524
332 524
3 2 66 0 0 12416 0 60 59 0 0 4
377 533
388 533
388 523
401 523
3 1 67 0 0 12416 0 61 59 0 0 4
382 497
389 497
389 505
401 505
1 2 39 0 0 0 0 68 70 0 0 4
615 383
537 383
537 433
554 433
0 1 68 0 0 4096 0 0 70 132 0 3
547 402
547 415
554 415
3 0 69 0 0 4096 0 74 0 0 128 3
446 412
475 412
475 411
2 1 69 0 0 8320 0 67 69 0 0 4
483 411
475 411
475 442
481 442
1 1 2 0 0 0 0 72 75 0 0 4
336 386
262 386
262 423
269 423
3 1 70 0 0 12416 0 70 71 0 0 4
599 424
605 424
605 433
615 433
3 2 71 0 0 4224 0 69 71 0 0 2
526 451
615 451
3 2 68 0 0 4224 0 67 68 0 0 3
532 402
615 402
615 401
2 1 72 0 0 4224 0 75 73 0 0 4
305 423
328 423
328 422
331 422
3 2 73 0 0 12416 0 73 74 0 0 4
376 431
387 431
387 421
400 421
3 1 74 0 0 12416 0 72 74 0 0 4
381 395
388 395
388 403
400 403
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
909 431 1002 453
919 438 991 454
9 Carry-Bit
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1115 558 1174 580
1124 566 1164 582
5 0-XOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1115 580 1166 602
1124 587 1156 603
4 1-OR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1113 600 1172 622
1122 608 1162 624
5 2-AND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1112 622 1171 644
1121 629 1161 645
5 3-NOT
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
