CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
40
13 Logic Switch~
5 1035 637 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-32 -4 -18 4
2 V6
-1031 -637 -1017 -629
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7168 0 0
2
5.8997e-315 5.34643e-315
0
13 Logic Switch~
5 1035 667 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-30 -5 -16 3
2 V7
-1035 -667 -1021 -659
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3171 0 0
2
5.8997e-315 5.32571e-315
0
13 Logic Switch~
5 1133 152 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-35 -3 -21 5
2 V8
-1129 -150 -1115 -142
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4139 0 0
2
5.8997e-315 5.30499e-315
0
13 Logic Switch~
5 1034 338 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-30 -5 -16 3
2 V9
-1027 -340 -1013 -332
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6435 0 0
2
5.8997e-315 5.26354e-315
0
13 Logic Switch~
5 1038 310 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-30 -3 -16 5
3 V10
-1028 -310 -1007 -302
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5283 0 0
2
5.8997e-315 0
0
13 Logic Switch~
5 157 614 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-32 -4 -18 4
2 V5
-239 -617 -225 -609
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6874 0 0
2
5.8997e-315 5.26354e-315
0
13 Logic Switch~
5 157 644 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-30 -5 -16 3
2 V4
-225 -643 -211 -635
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5305 0 0
2
5.8997e-315 0
0
13 Logic Switch~
5 255 129 0 1 11
0 22
0
0 0 21360 0
2 0V
-35 -3 -21 5
2 V1
-255 -129 -241 -121
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
34 0 0
2
5.8997e-315 5.34643e-315
0
13 Logic Switch~
5 149 318 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-30 -5 -16 3
2 V3
-237 -102 -223 -94
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
969 0 0
2
5.8997e-315 0
0
13 Logic Switch~
5 150 287 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-30 -3 -16 5
2 V2
-147 -287 -133 -279
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8402 0 0
2
5.8997e-315 0
0
8 2-In OR~
219 1262 466 0 3 22
0 5 4 12
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3751 0 0
2
5.8997e-315 0
0
9 2-In AND~
219 1229 847 0 3 22
0 3 2 10
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
4292 0 0
2
5.8997e-315 0
0
9 2-In NOR~
219 1407 735 0 3 22
0 8 9 7
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U7B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
6118 0 0
2
5.8997e-315 0
0
9 2-In NOR~
219 1218 768 0 3 22
0 2 2 9
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
34 0 0
2
5.8997e-315 0
0
9 2-In NOR~
219 1216 702 0 3 22
0 3 3 8
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U6D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
6357 0 0
2
5.8997e-315 0
0
9 2-In NOR~
219 1364 380 0 3 22
0 11 11 13
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U6C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
319 0 0
2
5.8997e-315 0
0
9 2-In NOR~
219 1185 381 0 3 22
0 5 4 11
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U6B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3976 0 0
2
5.8997e-315 0
0
9 2-In NOR~
219 1261 121 0 3 22
0 6 6 14
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
7634 0 0
2
5.8997e-315 0
0
14 Logic Display~
6 1528 843 0 1 2
10 10
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L7
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
523 0 0
2
5.8997e-315 5.4371e-315
0
14 Logic Display~
6 1527 731 0 1 2
10 7
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L8
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6748 0 0
2
5.8997e-315 5.42414e-315
0
14 Logic Display~
6 1415 184 0 1 2
10 15
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L9
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6901 0 0
2
5.8997e-315 5.41378e-315
0
9 Inverter~
13 1268 188 0 2 22
0 6 15
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
842 0 0
2
5.8997e-315 5.4086e-315
0
14 Logic Display~
6 1414 117 0 1 2
10 14
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L10
-8 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3277 0 0
2
5.8997e-315 5.39824e-315
0
14 Logic Display~
6 1469 462 0 1 2
10 12
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L11
-8 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4212 0 0
2
5.8997e-315 5.39306e-315
0
14 Logic Display~
6 1469 376 0 1 2
10 13
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L12
-8 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4720 0 0
2
5.8997e-315 5.36716e-315
0
14 Logic Display~
6 650 819 0 1 2
10 18
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L6
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5551 0 0
2
5.8997e-315 0
0
10 2-In NAND~
219 533 715 0 3 22
0 21 20 19
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
6986 0 0
2
5.8997e-315 0
0
8 2-In OR~
219 340 823 0 3 22
0 17 16 18
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
8745 0 0
2
5.8997e-315 0
0
10 2-In NAND~
219 347 746 0 3 22
0 16 16 20
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
9592 0 0
2
5.8997e-315 5.30499e-315
0
14 Logic Display~
6 651 711 0 1 2
10 19
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L5
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8748 0 0
2
5.8997e-315 5.26354e-315
0
10 2-In NAND~
219 347 679 0 3 22
0 17 17 21
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7168 0 0
2
5.8997e-315 0
0
14 Logic Display~
6 537 161 0 1 2
10 24
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
631 0 0
2
5.8997e-315 5.32571e-315
0
9 Inverter~
13 390 165 0 2 22
0 22 24
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
9466 0 0
2
5.8997e-315 5.30499e-315
0
10 2-In NAND~
219 394 99 0 3 22
0 22 22 23
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3266 0 0
2
5.8997e-315 5.26354e-315
0
14 Logic Display~
6 535 95 0 1 2
10 23
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7693 0 0
2
5.8997e-315 0
0
14 Logic Display~
6 591 439 0 1 2
10 25
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L4
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3723 0 0
2
5.8997e-315 0
0
10 2-In NAND~
219 315 356 0 3 22
0 28 27 26
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3440 0 0
2
5.8997e-315 0
0
9 2-In AND~
219 387 443 0 3 22
0 28 27 25
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
6263 0 0
2
5.8997e-315 0
0
14 Logic Display~
6 593 354 0 1 2
10 29
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L3
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4900 0 0
2
5.8997e-315 5.26354e-315
0
10 2-In NAND~
219 490 358 0 3 22
0 26 26 29
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
8783 0 0
2
5.8997e-315 0
0
46
0 0 2 0 0 4096 0 0 0 6 8 2
1125 768
1072 768
0 0 3 0 0 4096 0 0 0 7 9 2
1127 702
1047 702
2 0 4 0 0 4096 0 17 0 0 14 2
1172 390
1066 390
1 0 5 0 0 4096 0 17 0 0 15 2
1172 372
1047 372
1 0 6 0 0 8192 0 3 0 0 22 4
1145 152
1150 152
1150 121
1155 121
1 2 2 0 0 4096 0 14 14 0 0 4
1205 759
1125 759
1125 777
1205 777
1 2 3 0 0 0 0 15 15 0 0 4
1203 693
1127 693
1127 711
1203 711
1 2 2 0 0 8320 0 1 12 0 0 4
1047 637
1072 637
1072 856
1205 856
1 1 3 0 0 4224 0 2 12 0 0 3
1047 667
1047 838
1205 838
3 1 7 0 0 4224 0 13 20 0 0 2
1446 735
1511 735
3 1 8 0 0 4224 0 15 13 0 0 4
1255 702
1380 702
1380 726
1394 726
3 2 9 0 0 4224 0 14 13 0 0 4
1257 768
1380 768
1380 744
1394 744
3 1 10 0 0 4224 0 12 19 0 0 2
1250 847
1512 847
1 2 4 0 0 12416 0 5 11 0 0 4
1050 310
1066 310
1066 475
1249 475
1 1 5 0 0 12416 0 4 11 0 0 4
1046 338
1047 338
1047 457
1249 457
0 3 11 0 0 4096 0 0 17 19 0 2
1280 381
1224 381
3 1 12 0 0 4224 0 11 24 0 0 2
1295 466
1453 466
3 1 13 0 0 4224 0 16 25 0 0 2
1403 380
1453 380
1 2 11 0 0 4224 0 16 16 0 0 4
1351 371
1280 371
1280 389
1351 389
3 1 14 0 0 4224 0 18 23 0 0 2
1300 121
1398 121
1 1 6 0 0 4224 0 22 3 0 0 4
1253 188
1150 188
1150 152
1145 152
1 2 6 0 0 0 0 18 18 0 0 4
1248 112
1155 112
1155 130
1248 130
1 2 15 0 0 4224 0 21 22 0 0 2
1399 188
1289 188
0 0 16 0 0 4096 0 0 0 30 32 2
254 745
189 745
0 0 17 0 0 4096 0 0 0 31 33 2
251 679
169 679
3 1 18 0 0 4224 0 28 26 0 0 2
373 823
634 823
3 1 19 0 0 4224 0 27 30 0 0 2
560 715
635 715
2 3 20 0 0 12416 0 27 29 0 0 4
509 724
447 724
447 746
374 746
3 1 21 0 0 4224 0 31 27 0 0 4
374 679
448 679
448 706
509 706
1 2 16 0 0 4096 0 29 29 0 0 4
323 737
254 737
254 755
323 755
1 2 17 0 0 0 0 31 31 0 0 4
323 670
251 670
251 688
323 688
1 2 16 0 0 8320 0 6 28 0 0 4
169 614
189 614
189 832
327 832
1 1 17 0 0 4224 0 7 28 0 0 3
169 644
169 814
327 814
1 0 22 0 0 4096 0 8 0 0 35 2
267 129
290 129
1 0 22 0 0 4224 0 33 0 0 38 3
375 165
290 165
290 108
1 3 23 0 0 4224 0 35 34 0 0 2
519 99
421 99
1 2 24 0 0 4224 0 32 33 0 0 2
521 165
411 165
1 2 22 0 0 0 0 34 34 0 0 4
370 90
290 90
290 108
370 108
3 1 25 0 0 4224 0 38 36 0 0 2
408 443
575 443
0 3 26 0 0 4096 0 0 37 46 0 2
403 356
342 356
2 0 27 0 0 4096 0 37 0 0 43 2
291 365
183 365
1 0 28 0 0 4096 0 37 0 0 44 2
291 347
162 347
1 2 27 0 0 12416 0 10 38 0 0 4
162 287
183 287
183 452
363 452
1 1 28 0 0 12416 0 9 38 0 0 4
161 318
162 318
162 434
363 434
1 3 29 0 0 4224 0 39 40 0 0 2
577 358
517 358
1 2 26 0 0 4224 0 40 40 0 0 4
466 349
403 349
403 367
466 367
116
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
508 359 577 383
518 367 566 383
6 Pin- 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
402 360 471 384
412 368 460 384
6 Pin- 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
404 323 473 347
414 331 462 347
6 Pin- 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
79 302 124 326
89 310 113 326
3 A =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
79 273 124 297
89 281 113 297
3 B =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
222 324 291 348
232 332 280 348
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
222 358 291 382
232 366 280 382
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
332 360 401 384
342 368 390 384
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
239 407 308 431
249 415 297 431
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
239 446 308 470
249 454 297 470
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
409 441 478 465
419 449 467 465
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
191 408 220 432
201 416 209 432
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
191 445 220 469
201 453 209 469
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
188 319 217 343
198 327 206 343
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
188 358 217 382
198 366 206 382
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
349 326 386 350
359 334 375 350
2 AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
524 329 561 353
534 337 550 353
2 AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
441 415 478 439
451 423 467 439
2 AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
345 310 390 334
355 318 379 334
3 ___
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
275 479 424 503
285 487 413 503
16 NAND gate as AND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
300 64 369 88
310 72 358 88
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
298 103 367 127
308 111 356 127
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
416 92 485 116
426 100 474 116
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
298 158 367 182
308 166 356 182
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
417 158 486 182
427 166 475 182
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
325 137 354 161
335 145 343 161
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
422 70 451 94
432 78 440 94
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
426 142 455 166
436 150 444 166
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
418 55 455 79
428 63 444 79
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
422 127 459 151
432 135 448 151
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
313 83 342 107
323 91 331 107
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
182 113 227 137
192 121 216 137
3 A =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
316 191 465 215
326 199 454 215
16 NAND gate as NOT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
88 597 133 621
98 605 122 621
3 B =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
88 628 133 652
98 636 122 652
3 A =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
363 672 432 696
373 680 421 696
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
260 680 329 704
270 688 318 704
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
258 647 327 671
268 655 316 671
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
256 714 325 738
266 722 314 738
6 Pin- 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
256 748 325 772
266 756 314 772
6 Pin- 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
368 738 437 762
378 746 426 762
6 Pin- 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
443 682 512 706
453 690 501 706
6 Pin- 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
443 715 512 739
453 723 501 739
6 Pin-10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
557 710 626 734
567 718 615 734
6 Pin- 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
243 788 312 812
253 796 301 812
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
243 828 312 852
253 836 301 852
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
414 818 483 842
424 826 472 842
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
198 787 227 811
208 795 216 811
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
199 828 228 852
209 836 217 852
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
204 655 233 679
214 663 222 679
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
203 721 232 745
213 729 221 745
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
383 638 420 662
393 646 409 662
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
387 653 416 677
397 661 405 677
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
383 707 420 731
393 715 409 731
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
388 721 413 745
396 729 404 745
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
559 686 620 710
569 694 609 710
5 A + B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
422 792 483 816
432 800 472 816
5 A + B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
277 875 418 899
287 883 407 899
15 NAND gate as OR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
966 322 1011 346
976 330 1000 346
3 A =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
965 295 1010 319
975 303 999 319
3 B =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1117 430 1186 454
1127 438 1175 454
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1117 469 1186 493
1127 477 1175 493
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1316 464 1385 488
1326 472 1374 488
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1069 431 1098 455
1079 439 1087 455
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1069 468 1098 492
1079 476 1087 492
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1066 342 1095 366
1076 350 1084 366
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1066 381 1095 405
1076 389 1084 405
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1451 709 1488 733
1461 717 1477 733
2 AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1226 339 1271 363
1236 347 1260 363
3 ___
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1176 181 1245 205
1186 189 1234 205
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1295 181 1364 205
1305 189 1353 205
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1203 160 1232 184
1213 168 1221 184
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1300 93 1329 117
1310 101 1318 117
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1304 165 1333 189
1314 173 1322 189
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1296 78 1333 102
1306 86 1322 102
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1300 150 1337 174
1310 158 1326 174
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1191 106 1220 130
1201 114 1209 130
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1060 136 1105 160
1070 144 1094 160
3 A =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
966 620 1011 644
976 628 1000 644
3 B =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
966 651 1011 675
976 659 1000 675
3 A =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1121 811 1190 835
1131 819 1179 835
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1121 851 1190 875
1131 859 1179 875
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1292 841 1361 865
1302 849 1350 865
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1076 810 1105 834
1086 818 1094 834
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1077 851 1106 875
1087 859 1095 875
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1082 678 1111 702
1092 686 1100 702
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1081 744 1110 768
1091 752 1099 768
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1261 661 1298 685
1271 669 1287 685
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1265 676 1294 700
1275 684 1283 700
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1261 730 1298 754
1271 738 1287 754
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1266 744 1291 768
1274 752 1282 768
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1178 87 1245 109
1187 95 1235 111
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1176 126 1243 148
1185 134 1233 150
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1294 115 1361 137
1303 123 1351 139
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
1194 214 1333 236
1203 221 1323 237
15 NOR gate as NOT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1100 347 1167 369
1109 355 1157 371
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1099 385 1166 407
1108 393 1156 409
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1210 383 1277 405
1219 390 1267 406
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1282 346 1349 368
1291 354 1339 370
6 Pin- 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1284 383 1351 405
1293 390 1341 406
6 Pin- 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1394 376 1461 398
1403 384 1451 400
6 Pin- 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1227 357 1270 379
1236 364 1260 380
3 A+B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1406 355 1449 377
1415 362 1439 378
3 A+B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1322 441 1383 465
1332 449 1372 465
5 A + B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1310 818 1347 842
1320 826 1336 842
2 AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1136 670 1203 692
1145 677 1193 693
6 Pin- 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1141 703 1208 725
1150 710 1198 726
6 Pin- 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1241 695 1308 717
1250 703 1298 719
6 Pin- 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1134 737 1201 759
1143 745 1191 761
6 Pin- 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1134 771 1201 793
1143 778 1191 794
6 Pin- 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1246 761 1313 783
1255 768 1303 784
6 Pin- 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1316 696 1383 718
1325 704 1373 720
6 Pin- 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1324 742 1383 764
1333 749 1373 765
5 Pin-9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1440 733 1515 755
1449 740 1505 756
7 Pin- 10
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 14
1153 502 1298 527
1162 509 1288 526
14 NOR gate as OR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
1155 898 1296 920
1165 905 1285 921
15 NOR gate as AND
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
