CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
1090 790 30 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
176 502 1364 707
9437202 0
0
6 Title:
5 Name:
0
0
0
159
13 Logic Switch~
5 1243 1205 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 E1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3947 0 0
2
5.89976e-315 0
0
13 Logic Switch~
5 1120 1050 0 10 11
0 71 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 F
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5715 0 0
2
5.89976e-315 5.3568e-315
0
13 Logic Switch~
5 1209 1050 0 10 11
0 68 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 C
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5703 0 0
2
5.89976e-315 5.34643e-315
0
13 Logic Switch~
5 1233 1049 0 1 11
0 69
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3511 0 0
2
5.89976e-315 5.32571e-315
0
13 Logic Switch~
5 1259 1048 0 10 11
0 70 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9901 0 0
2
5.89976e-315 5.30499e-315
0
13 Logic Switch~
5 1178 1051 0 10 11
0 73 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 D
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9115 0 0
2
5.89976e-315 5.26354e-315
0
13 Logic Switch~
5 1146 1052 0 1 11
0 72
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 E
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5545 0 0
2
5.89976e-315 0
0
13 Logic Switch~
5 1784 639 0 1 11
0 118
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9700 0 0
2
5.89976e-315 0
0
13 Logic Switch~
5 1749 639 0 10 11
0 119 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3905 0 0
2
5.89976e-315 0
0
13 Logic Switch~
5 1030 596 0 10 11
0 120 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 E
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
976 0 0
2
5.89976e-315 0
0
13 Logic Switch~
5 1062 595 0 10 11
0 121 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 D
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3676 0 0
2
5.89976e-315 0
0
13 Logic Switch~
5 1143 592 0 1 11
0 124
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6137 0 0
2
5.89976e-315 5.30499e-315
0
13 Logic Switch~
5 1117 593 0 10 11
0 123 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3458 0 0
2
5.89976e-315 5.26354e-315
0
13 Logic Switch~
5 1093 594 0 10 11
0 122 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 C
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8160 0 0
2
5.89976e-315 0
0
13 Logic Switch~
5 119 794 0 1 11
0 128
0
0 0 21360 0
2 0V
-27 -6 -13 2
2 V8
-40 43 -26 51
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8874 0 0
2
44262.9 0
0
13 Logic Switch~
5 119 766 0 10 11
0 129 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-32 0 -18 8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3791 0 0
2
44262.9 1
0
13 Logic Switch~
5 120 578 0 1 11
0 125
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 C
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9555 0 0
2
44262.9 2
0
13 Logic Switch~
5 150 579 0 10 11
0 126 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3215 0 0
2
44262.9 3
0
13 Logic Switch~
5 179 582 0 1 11
0 127
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7300 0 0
2
44262.9 4
0
13 Logic Switch~
5 475 80 0 10 11
0 141 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
587 58 601 66
2 V3
536 -3 550 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3165 0 0
2
44262.9 5
0
13 Logic Switch~
5 78 116 0 10 11
0 140 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-36 -7 -22 1
2 V2
-67 -6 -53 2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7874 0 0
2
44262.9 6
0
13 Logic Switch~
5 79 61 0 10 11
0 139 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-34 -7 -20 1
2 V1
-64 -10 -50 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3280 0 0
2
44262.9 7
0
14 Logic Display~
6 1289 967 0 1 2
10 58
0
0 0 53872 90
6 100MEG
3 -16 45 -8
4 L108
1265 -81 1293 -73
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3122 0 0
2
5.89976e-315 5.36716e-315
0
14 Logic Display~
6 1288 945 0 1 2
10 57
0
0 0 53872 90
6 100MEG
3 -16 45 -8
4 L107
1149 -100 1177 -92
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6242 0 0
2
5.89976e-315 5.3568e-315
0
14 Logic Display~
6 1288 922 0 1 2
10 56
0
0 0 53872 90
6 100MEG
3 -16 45 -8
4 L106
1198 47 1226 55
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8862 0 0
2
5.89976e-315 5.34643e-315
0
14 Logic Display~
6 1287 899 0 1 2
10 55
0
0 0 53872 90
6 100MEG
3 -16 45 -8
4 L105
1267 118 1295 126
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3202 0 0
2
5.89976e-315 5.32571e-315
0
14 Logic Display~
6 1287 879 0 1 2
10 54
0
0 0 53872 90
6 100MEG
3 -16 45 -8
4 L104
1247 59 1275 67
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5657 0 0
2
5.89976e-315 5.30499e-315
0
14 Logic Display~
6 1284 837 0 1 2
10 52
0
0 0 53872 90
6 100MEG
3 -16 45 -8
4 L103
1250 7 1278 15
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3554 0 0
2
5.89976e-315 5.26354e-315
0
14 Logic Display~
6 1284 857 0 1 2
10 53
0
0 0 53872 90
6 100MEG
3 -16 45 -8
4 L102
1168 165 1196 173
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4316 0 0
2
5.89976e-315 0
0
14 Logic Display~
6 1388 966 0 1 2
10 51
0
0 0 53872 90
6 100MEG
3 -16 45 -8
4 L101
1265 -81 1293 -73
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3739 0 0
2
5.89976e-315 5.36716e-315
0
14 Logic Display~
6 1387 944 0 1 2
10 50
0
0 0 53872 90
6 100MEG
3 -16 45 -8
4 L100
1149 -100 1177 -92
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7606 0 0
2
5.89976e-315 5.3568e-315
0
14 Logic Display~
6 1387 921 0 1 2
10 49
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L99
1201 47 1222 55
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3741 0 0
2
5.89976e-315 5.34643e-315
0
14 Logic Display~
6 1386 898 0 1 2
10 48
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L98
1270 118 1291 126
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
369 0 0
2
5.89976e-315 5.32571e-315
0
14 Logic Display~
6 1386 878 0 1 2
10 47
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L97
1250 59 1271 67
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8773 0 0
2
5.89976e-315 5.30499e-315
0
14 Logic Display~
6 1383 836 0 1 2
10 45
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L96
1253 7 1274 15
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7981 0 0
2
5.89976e-315 5.26354e-315
0
14 Logic Display~
6 1383 856 0 1 2
10 46
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L95
1171 165 1192 173
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4205 0 0
2
5.89976e-315 0
0
14 Logic Display~
6 1483 970 0 1 2
10 44
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L94
1268 -81 1289 -73
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3375 0 0
2
5.89976e-315 5.36716e-315
0
14 Logic Display~
6 1482 948 0 1 2
10 43
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L93
1152 -100 1173 -92
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
719 0 0
2
5.89976e-315 5.3568e-315
0
14 Logic Display~
6 1482 925 0 1 2
10 42
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L92
1201 47 1222 55
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3749 0 0
2
5.89976e-315 5.34643e-315
0
14 Logic Display~
6 1481 902 0 1 2
10 41
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L91
1270 118 1291 126
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3871 0 0
2
5.89976e-315 5.32571e-315
0
14 Logic Display~
6 1481 882 0 1 2
10 40
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L90
1250 59 1271 67
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4393 0 0
2
5.89976e-315 5.30499e-315
0
14 Logic Display~
6 1478 840 0 1 2
10 38
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L89
1253 7 1274 15
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6229 0 0
2
5.89976e-315 5.26354e-315
0
14 Logic Display~
6 1478 860 0 1 2
10 39
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L88
1171 165 1192 173
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3757 0 0
2
5.89976e-315 0
0
14 Logic Display~
6 1572 858 0 1 2
10 32
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L87
1171 165 1192 173
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
352 0 0
2
5.89976e-315 5.36716e-315
0
14 Logic Display~
6 1572 838 0 1 2
10 31
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L86
1253 7 1274 15
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3372 0 0
2
5.89976e-315 5.3568e-315
0
14 Logic Display~
6 1575 880 0 1 2
10 33
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L85
1250 59 1271 67
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4911 0 0
2
5.89976e-315 5.34643e-315
0
14 Logic Display~
6 1575 900 0 1 2
10 34
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L84
1270 118 1291 126
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7574 0 0
2
5.89976e-315 5.32571e-315
0
14 Logic Display~
6 1576 923 0 1 2
10 35
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L83
1201 47 1222 55
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6601 0 0
2
5.89976e-315 5.30499e-315
0
14 Logic Display~
6 1576 946 0 1 2
10 36
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L82
1152 -100 1173 -92
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8531 0 0
2
5.89976e-315 5.26354e-315
0
14 Logic Display~
6 1577 968 0 1 2
10 37
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L81
1268 -81 1289 -73
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6532 0 0
2
5.89976e-315 0
0
14 Logic Display~
6 1667 856 0 1 2
10 25
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L80
1178 102 1199 110
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3621 0 0
2
5.89976e-315 5.36716e-315
0
14 Logic Display~
6 1667 836 0 1 2
10 24
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L79
1018 34 1039 42
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5174 0 0
2
5.89976e-315 5.3568e-315
0
14 Logic Display~
6 1670 878 0 1 2
10 26
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L78
1092 -32 1113 -24
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5452 0 0
2
5.89976e-315 5.34643e-315
0
14 Logic Display~
6 1670 898 0 1 2
10 27
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L77
1175 118 1196 126
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3626 0 0
2
5.89976e-315 5.32571e-315
0
14 Logic Display~
6 1671 921 0 1 2
10 28
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L76
1174 101 1195 109
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3806 0 0
2
5.89976e-315 5.30499e-315
0
14 Logic Display~
6 1671 944 0 1 2
10 29
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L75
1174 9 1195 17
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3389 0 0
2
5.89976e-315 5.26354e-315
0
14 Logic Display~
6 1672 966 0 1 2
10 30
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L74
972 -147 993 -139
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9156 0 0
2
5.89976e-315 0
0
14 Logic Display~
6 1764 863 0 1 2
10 18
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L73
471 119 492 127
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5810 0 0
2
5.89976e-315 5.36716e-315
0
14 Logic Display~
6 1764 843 0 1 2
10 17
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L72
454 54 475 62
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8260 0 0
2
5.89976e-315 5.3568e-315
0
14 Logic Display~
6 1767 885 0 1 2
10 19
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L71
454 54 475 62
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7286 0 0
2
5.89976e-315 5.34643e-315
0
14 Logic Display~
6 1767 905 0 1 2
10 20
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L70
471 119 492 127
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3689 0 0
2
5.89976e-315 5.32571e-315
0
14 Logic Display~
6 1768 928 0 1 2
10 21
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L69
481 101 502 109
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4485 0 0
2
5.89976e-315 5.30499e-315
0
14 Logic Display~
6 1768 951 0 1 2
10 22
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L68
449 26 470 34
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4370 0 0
2
5.89976e-315 5.26354e-315
0
14 Logic Display~
6 1769 973 0 1 2
10 23
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L67
493 -28 514 -20
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7483 0 0
2
5.89976e-315 0
0
14 Logic Display~
6 1868 974 0 1 2
10 16
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L66
493 -28 514 -20
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4214 0 0
2
5.89976e-315 5.36716e-315
0
14 Logic Display~
6 1867 952 0 1 2
10 15
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L65
449 26 470 34
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9254 0 0
2
5.89976e-315 5.3568e-315
0
14 Logic Display~
6 1867 929 0 1 2
10 14
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L64
481 101 502 109
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7515 0 0
2
5.89976e-315 5.34643e-315
0
14 Logic Display~
6 1866 906 0 1 2
10 13
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L61
471 119 492 127
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9241 0 0
2
5.89976e-315 5.32571e-315
0
14 Logic Display~
6 1866 886 0 1 2
10 12
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L60
454 54 475 62
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3783 0 0
2
5.89976e-315 5.30499e-315
0
14 Logic Display~
6 1863 844 0 1 2
10 10
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L59
454 54 475 62
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5226 0 0
2
5.89976e-315 5.26354e-315
0
14 Logic Display~
6 1863 864 0 1 2
10 11
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L58
471 119 492 127
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6496 0 0
2
5.89976e-315 0
0
14 Logic Display~
6 1957 854 0 1 2
10 4
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L63
471 119 492 127
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6819 0 0
2
5.89976e-315 5.26354e-315
0
14 Logic Display~
6 1957 834 0 1 2
10 3
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L62
454 54 475 62
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6832 0 0
2
5.89976e-315 0
0
14 Logic Display~
6 1960 876 0 1 2
10 5
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L57
454 54 475 62
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7222 0 0
2
5.89976e-315 5.26354e-315
0
14 Logic Display~
6 1960 896 0 1 2
10 6
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L56
471 119 492 127
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4676 0 0
2
5.89976e-315 0
0
14 Logic Display~
6 1961 919 0 1 2
10 7
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L55
481 101 502 109
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9334 0 0
2
5.89976e-315 5.26354e-315
0
14 Logic Display~
6 1961 942 0 1 2
10 8
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L54
449 26 470 34
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4758 0 0
2
5.89976e-315 0
0
14 Logic Display~
6 1964 988 0 1 2
10 59
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L53
473 2 494 10
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6695 0 0
2
5.89976e-315 5.38788e-315
0
14 Logic Display~
6 1869 992 0 1 2
10 60
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L52
586 77 607 85
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8212 0 0
2
5.89976e-315 5.37752e-315
0
14 Logic Display~
6 1770 995 0 1 2
10 61
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L51
507 90 528 98
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3922 0 0
2
5.89976e-315 5.36716e-315
0
14 Logic Display~
6 1671 992 0 1 2
10 62
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L50
775 126 796 134
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7610 0 0
2
5.89976e-315 5.3568e-315
0
14 Logic Display~
6 1578 993 0 1 2
10 63
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L49
1267 82 1288 90
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6131 0 0
2
5.89976e-315 5.34643e-315
0
14 Logic Display~
6 1485 994 0 1 2
10 64
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L48
999 -187 1020 -179
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7187 0 0
2
5.89976e-315 5.32571e-315
0
14 Logic Display~
6 1386 995 0 1 2
10 65
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L47
1475 -121 1496 -113
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9198 0 0
2
5.89976e-315 5.30499e-315
0
14 Logic Display~
6 1291 990 0 1 2
10 66
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L46
1574 65 1595 73
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9468 0 0
2
5.89976e-315 5.26354e-315
0
14 Logic Display~
6 1962 964 0 1 2
10 9
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 L45
493 -28 514 -20
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5160 0 0
2
5.89976e-315 0
0
9 Inverter~
13 1338 1228 0 2 22
0 2 67
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 4 0
1 U
7647 0 0
2
5.89976e-315 0
0
7 74LS138
19 1697 1213 0 14 29
0 71 72 73 2 67 67 81 80 79
78 77 76 75 74
0
0 0 5104 90
6 74F138
-22 -8 20 0
3 U19
-761 -358 -740 -350
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
7210 0 0
2
5.89976e-315 0
0
7 74LS138
19 1715 1067 0 14 29
0 68 69 70 2 77 77 62 30 29
28 27 26 25 24
0
0 0 5104 90
6 74F138
-14 -9 28 -1
3 U18
-767 -208 -746 -200
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
7128 0 0
2
5.89976e-315 5.32571e-315
0
7 74LS138
19 1811 1068 0 14 29
0 68 69 70 2 76 76 61 23 22
21 20 19 18 17
0
0 0 5104 90
6 74F138
-22 -8 20 0
3 U17
-853 -220 -832 -212
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
5367 0 0
2
5.89976e-315 5.30499e-315
0
7 74LS138
19 2002 1068 0 14 29
0 68 69 70 2 74 74 59 9 8
7 6 5 4 3
0
0 0 5104 90
6 74F138
-20 -7 22 1
3 U16
-1089 -216 -1068 -208
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
7140 0 0
2
5.89976e-315 5.26354e-315
0
7 74LS138
19 1907 1068 0 14 29
0 68 69 70 2 75 75 60 16 15
14 13 12 11 10
0
0 0 5104 90
6 74F138
-17 -9 25 -1
3 U15
-952 -194 -931 -186
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
4903 0 0
2
5.89976e-315 0
0
7 74LS138
19 1331 1066 0 14 29
0 68 69 70 2 81 81 66 58 57
56 55 54 53 52
0
0 0 5104 90
6 74F138
-14 -9 28 -1
3 U14
-350 -169 -329 -161
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
3690 0 0
2
5.89976e-315 5.32571e-315
0
7 74LS138
19 1427 1066 0 14 29
0 68 69 70 2 80 80 65 51 50
49 48 47 46 45
0
0 0 5104 90
6 74F138
-22 -8 20 0
3 U13
-499 -180 -478 -172
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
8598 0 0
2
5.89976e-315 5.30499e-315
0
7 74LS138
19 1619 1067 0 14 29
0 68 69 70 2 78 78 63 37 36
35 34 33 32 31
0
0 0 5104 90
6 74F138
-20 -7 22 1
3 U12
-605 -230 -584 -222
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
5737 0 0
2
5.89976e-315 5.26354e-315
0
7 74LS138
19 1523 1067 0 14 29
0 68 69 70 2 79 79 64 44 43
42 41 40 39 38
0
0 0 5104 90
6 74F138
-17 -9 25 -1
3 U11
-503 -190 -482 -182
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
3882 0 0
2
5.89976e-315 0
0
14 Logic Display~
6 1504 430 0 1 2
10 98
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3440 0 0
2
5.89976e-315 5.46818e-315
0
14 Logic Display~
6 1479 431 0 1 2
10 99
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5176 0 0
2
5.89976e-315 5.46559e-315
0
14 Logic Display~
6 1452 430 0 1 2
10 100
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9582 0 0
2
5.89976e-315 5.463e-315
0
14 Logic Display~
6 1427 430 0 1 2
10 101
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9862 0 0
2
5.89976e-315 5.46041e-315
0
14 Logic Display~
6 1403 432 0 1 2
10 102
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5432 0 0
2
5.89976e-315 5.45782e-315
0
14 Logic Display~
6 1379 431 0 1 2
10 103
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L18
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3602 0 0
2
5.89976e-315 5.45523e-315
0
14 Logic Display~
6 1353 432 0 1 2
10 104
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4714 0 0
2
5.89976e-315 5.45264e-315
0
14 Logic Display~
6 1330 432 0 1 2
10 105
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L20
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3834 0 0
2
5.89976e-315 5.45005e-315
0
14 Logic Display~
6 1304 433 0 1 2
10 106
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L21
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3577 0 0
2
5.89976e-315 5.44746e-315
0
14 Logic Display~
6 1279 434 0 1 2
10 107
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L22
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7571 0 0
2
5.89976e-315 5.44487e-315
0
14 Logic Display~
6 1253 435 0 1 2
10 108
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L23
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
311 0 0
2
5.89976e-315 5.44228e-315
0
14 Logic Display~
6 1227 435 0 1 2
10 109
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L24
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5524 0 0
2
5.89976e-315 5.43969e-315
0
14 Logic Display~
6 1203 435 0 1 2
10 110
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L25
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6424 0 0
2
5.89976e-315 5.4371e-315
0
14 Logic Display~
6 1178 436 0 1 2
10 111
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L26
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8878 0 0
2
5.89976e-315 5.43451e-315
0
14 Logic Display~
6 1153 436 0 1 2
10 112
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L27
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3615 0 0
2
5.89976e-315 5.43192e-315
0
14 Logic Display~
6 1130 437 0 1 2
10 113
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L28
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7948 0 0
2
5.89976e-315 5.42933e-315
0
14 Logic Display~
6 1523 430 0 1 2
10 97
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L29
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
447 0 0
2
5.89976e-315 5.42414e-315
0
14 Logic Display~
6 1546 429 0 1 2
10 96
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L30
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4827 0 0
2
5.89976e-315 5.41896e-315
0
14 Logic Display~
6 1571 429 0 1 2
10 95
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L31
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3675 0 0
2
5.89976e-315 5.41378e-315
0
14 Logic Display~
6 1596 428 0 1 2
10 94
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L32
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7278 0 0
2
5.89976e-315 5.4086e-315
0
14 Logic Display~
6 1620 428 0 1 2
10 93
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L33
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
926 0 0
2
5.89976e-315 5.40342e-315
0
14 Logic Display~
6 1646 428 0 1 2
10 92
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L34
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6747 0 0
2
5.89976e-315 5.39824e-315
0
14 Logic Display~
6 1672 427 0 1 2
10 91
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L35
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5177 0 0
2
5.89976e-315 5.39306e-315
0
14 Logic Display~
6 1697 426 0 1 2
10 90
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L36
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5594 0 0
2
5.89976e-315 5.38788e-315
0
14 Logic Display~
6 1723 425 0 1 2
10 89
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L37
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9933 0 0
2
5.89976e-315 5.37752e-315
0
14 Logic Display~
6 1746 425 0 1 2
10 88
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L38
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8987 0 0
2
5.89976e-315 5.36716e-315
0
14 Logic Display~
6 1772 424 0 1 2
10 87
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L39
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3275 0 0
2
5.89976e-315 5.3568e-315
0
14 Logic Display~
6 1796 425 0 1 2
10 86
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L40
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3551 0 0
2
5.89976e-315 5.34643e-315
0
14 Logic Display~
6 1820 423 0 1 2
10 85
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L41
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9522 0 0
2
5.89976e-315 5.32571e-315
0
14 Logic Display~
6 1845 423 0 1 2
10 84
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L42
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3443 0 0
2
5.89976e-315 5.30499e-315
0
14 Logic Display~
6 1872 424 0 1 2
10 83
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L43
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3935 0 0
2
5.89976e-315 5.26354e-315
0
14 Logic Display~
6 1897 423 0 1 2
10 82
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L44
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4532 0 0
2
5.89976e-315 0
0
7 74LS138
19 1461 723 0 14 29
0 118 120 121 119 118 118 154 155 156
157 114 115 116 117
0
0 0 5104 90
6 74F138
-14 -9 28 -1
3 U10
-125 -18 -104 -10
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 512 1 0 0 0
1 U
7600 0 0
2
5.89976e-315 0
0
7 74LS138
19 1524 585 0 14 29
0 122 123 124 119 116 116 97 96 95
94 93 92 91 90
0
0 0 5104 90
6 74F138
-17 -9 25 -1
2 U9
-500 -190 -486 -182
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
6952 0 0
2
5.89976e-315 5.43192e-315
0
7 74LS138
19 1624 584 0 14 29
0 122 123 124 119 117 117 89 88 87
86 85 84 83 82
0
0 0 5104 90
6 74F138
-20 -7 22 1
2 U8
-602 -230 -588 -222
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
3663 0 0
2
5.89976e-315 5.42933e-315
0
7 74LS138
19 1390 587 0 14 29
0 122 123 124 119 115 115 105 104 103
102 101 100 99 98
0
0 0 5104 90
6 74F138
-22 -8 20 0
2 U7
-496 -180 -482 -172
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
9511 0 0
2
5.89976e-315 0
0
7 74LS138
19 1275 587 0 14 29
0 122 123 124 119 114 114 113 112 111
110 109 108 107 106
0
0 0 5104 90
6 74F138
-14 -9 28 -1
2 U6
-347 -169 -333 -161
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
4625 0 0
2
5.89976e-315 0
0
14 Logic Display~
6 762 607 0 1 2
10 137
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6215 0 0
2
44262.9 8
0
14 Logic Display~
6 736 607 0 1 2
10 136
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4535 0 0
2
44262.9 9
0
14 Logic Display~
6 707 609 0 1 2
10 135
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3611 0 0
2
44262.9 10
0
14 Logic Display~
6 685 611 0 1 2
10 134
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9183 0 0
2
44262.9 11
0
14 Logic Display~
6 661 611 0 1 2
10 133
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3593 0 0
2
44262.9 12
0
14 Logic Display~
6 636 612 0 1 2
10 132
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4142 0 0
2
44262.9 13
0
14 Logic Display~
6 611 612 0 1 2
10 131
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9564 0 0
2
44262.9 14
0
14 Logic Display~
6 588 613 0 1 2
10 130
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7772 0 0
2
44262.9 15
0
7 74LS138
19 474 692 0 14 29
0 125 126 127 129 128 128 130 131 132
133 134 135 136 137
0
0 0 5104 0
6 74F138
-21 -61 21 -53
2 U5
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
3826 0 0
2
44262.9 16
0
9 Inverter~
13 170 223 0 2 22
0 139 138
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
9216 0 0
2
44262.9 17
0
9 Inverter~
13 461 345 0 2 22
0 138 146
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
770 0 0
2
44262.9 18
0
9 Inverter~
13 468 237 0 2 22
0 139 147
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
6894 0 0
2
44262.9 19
0
9 Inverter~
13 472 150 0 2 22
0 140 148
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
3840 0 0
2
44262.9 20
0
9 Inverter~
13 472 53 0 2 22
0 139 149
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
6568 0 0
2
44262.9 21
0
14 Logic Display~
6 780 324 0 1 2
10 142
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
656 0 0
2
44262.9 22
0
14 Logic Display~
6 784 231 0 1 2
10 143
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5430 0 0
2
44262.9 23
0
14 Logic Display~
6 779 138 0 1 2
10 144
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6853 0 0
2
44262.9 24
0
14 Logic Display~
6 779 47 0 1 2
10 145
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3322 0 0
2
44262.9 25
0
9 Inverter~
13 460 318 0 2 22
0 138 150
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
9236 0 0
2
44262.9 26
0
9 Inverter~
13 468 212 0 2 22
0 139 151
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
8728 0 0
2
44262.9 27
0
9 Inverter~
13 472 120 0 2 22
0 140 152
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
4790 0 0
2
44262.9 28
0
9 Inverter~
13 473 27 0 2 22
0 140 153
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3447 0 0
2
44262.9 29
0
5 4073~
219 619 354 0 4 22
0 150 146 140 142
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
4769 0 0
2
44262.9 30
0
5 4073~
219 615 251 0 4 22
0 151 147 140 143
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 1 0
1 U
3989 0 0
2
44262.9 31
0
5 4073~
219 614 162 0 4 22
0 152 148 139 144
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 1 0
1 U
3188 0 0
2
44262.9 32
0
5 4073~
219 608 70 0 4 22
0 153 149 141 145
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 1 0
1 U
7596 0 0
2
44262.9 33
0
220
4 0 2 0 0 12288 0 89 0 0 78 4
1736 1096
1736 1140
1764 1140
1764 1271
1 14 3 0 0 8320 0 73 91 0 0 3
1972 837
2041 837
2041 1027
1 13 4 0 0 8320 0 72 91 0 0 3
1972 857
2032 857
2032 1027
1 12 5 0 0 8320 0 74 91 0 0 3
1975 879
2023 879
2023 1027
1 11 6 0 0 8320 0 75 91 0 0 3
1975 899
2014 899
2014 1027
1 10 7 0 0 8320 0 76 91 0 0 3
1976 922
2005 922
2005 1027
1 9 8 0 0 8320 0 77 91 0 0 3
1976 945
1996 945
1996 1027
1 8 9 0 0 8320 0 86 91 0 0 3
1977 967
1987 967
1987 1027
1 14 10 0 0 8320 0 70 92 0 0 5
1878 847
1934 847
1934 1019
1946 1019
1946 1027
1 13 11 0 0 8320 0 71 92 0 0 3
1878 867
1937 867
1937 1027
1 12 12 0 0 8320 0 69 92 0 0 3
1881 889
1928 889
1928 1027
1 11 13 0 0 8320 0 68 92 0 0 3
1881 909
1919 909
1919 1027
1 10 14 0 0 8320 0 67 92 0 0 3
1882 932
1910 932
1910 1027
1 9 15 0 0 8320 0 66 92 0 0 3
1882 955
1901 955
1901 1027
1 8 16 0 0 8320 0 65 92 0 0 3
1883 977
1892 977
1892 1027
1 14 17 0 0 8320 0 59 90 0 0 5
1779 846
1845 846
1845 1019
1850 1019
1850 1027
1 13 18 0 0 8320 0 58 90 0 0 3
1779 866
1841 866
1841 1027
1 12 19 0 0 8320 0 60 90 0 0 3
1782 888
1832 888
1832 1027
1 11 20 0 0 8320 0 61 90 0 0 3
1782 908
1823 908
1823 1027
1 10 21 0 0 8320 0 62 90 0 0 3
1783 931
1814 931
1814 1027
1 9 22 0 0 8320 0 63 90 0 0 3
1783 954
1805 954
1805 1027
1 8 23 0 0 8320 0 64 90 0 0 3
1784 976
1796 976
1796 1027
1 14 24 0 0 8320 0 52 89 0 0 5
1682 839
1741 839
1741 1018
1754 1018
1754 1026
1 13 25 0 0 8320 0 51 89 0 0 3
1682 859
1745 859
1745 1026
1 12 26 0 0 8320 0 53 89 0 0 3
1685 881
1736 881
1736 1026
1 11 27 0 0 8320 0 54 89 0 0 3
1685 901
1727 901
1727 1026
1 10 28 0 0 8320 0 55 89 0 0 3
1686 924
1718 924
1718 1026
1 9 29 0 0 8320 0 56 89 0 0 3
1686 947
1709 947
1709 1026
1 8 30 0 0 8320 0 57 89 0 0 3
1687 969
1700 969
1700 1026
1 14 31 0 0 8320 0 45 95 0 0 5
1587 841
1644 841
1644 1018
1658 1018
1658 1026
1 13 32 0 0 8320 0 44 95 0 0 3
1587 861
1649 861
1649 1026
1 12 33 0 0 8320 0 46 95 0 0 3
1590 883
1640 883
1640 1026
1 11 34 0 0 8320 0 47 95 0 0 3
1590 903
1631 903
1631 1026
1 10 35 0 0 8320 0 48 95 0 0 3
1591 926
1622 926
1622 1026
1 9 36 0 0 8320 0 49 95 0 0 3
1591 949
1613 949
1613 1026
1 8 37 0 0 8320 0 50 95 0 0 3
1592 971
1604 971
1604 1026
1 14 38 0 0 8320 0 42 96 0 0 5
1493 843
1549 843
1549 1018
1562 1018
1562 1026
1 13 39 0 0 8320 0 43 96 0 0 3
1493 863
1553 863
1553 1026
1 12 40 0 0 8320 0 41 96 0 0 3
1496 885
1544 885
1544 1026
1 11 41 0 0 8320 0 40 96 0 0 3
1496 905
1535 905
1535 1026
1 10 42 0 0 8320 0 39 96 0 0 3
1497 928
1526 928
1526 1026
1 9 43 0 0 8320 0 38 96 0 0 3
1497 951
1517 951
1517 1026
1 8 44 0 0 8320 0 37 96 0 0 3
1498 973
1508 973
1508 1026
1 14 45 0 0 8320 0 35 94 0 0 5
1398 839
1460 839
1460 1017
1466 1017
1466 1025
1 13 46 0 0 8320 0 36 94 0 0 3
1398 859
1457 859
1457 1025
1 12 47 0 0 8320 0 34 94 0 0 3
1401 881
1448 881
1448 1025
1 11 48 0 0 8320 0 33 94 0 0 3
1401 901
1439 901
1439 1025
1 10 49 0 0 8320 0 32 94 0 0 3
1402 924
1430 924
1430 1025
1 9 50 0 0 8320 0 31 94 0 0 3
1402 947
1421 947
1421 1025
1 8 51 0 0 8320 0 30 94 0 0 3
1403 969
1412 969
1412 1025
1 14 52 0 0 8320 0 28 93 0 0 5
1299 840
1365 840
1365 1017
1370 1017
1370 1025
1 13 53 0 0 8320 0 29 93 0 0 3
1299 860
1361 860
1361 1025
1 12 54 0 0 8320 0 27 93 0 0 3
1302 882
1352 882
1352 1025
1 11 55 0 0 8320 0 26 93 0 0 3
1302 902
1343 902
1343 1025
1 10 56 0 0 8320 0 25 93 0 0 3
1303 925
1334 925
1334 1025
1 9 57 0 0 8320 0 24 93 0 0 3
1303 948
1325 948
1325 1025
1 8 58 0 0 8320 0 23 93 0 0 3
1304 970
1316 970
1316 1025
1 7 59 0 0 8320 0 78 91 0 0 3
1979 991
1978 991
1978 1027
1 7 60 0 0 8320 0 79 92 0 0 3
1884 995
1883 995
1883 1027
1 7 61 0 0 8320 0 80 90 0 0 3
1785 998
1787 998
1787 1027
1 7 62 0 0 8320 0 81 89 0 0 3
1686 995
1691 995
1691 1026
1 7 63 0 0 8320 0 82 95 0 0 3
1593 996
1595 996
1595 1026
1 7 64 0 0 8320 0 83 96 0 0 3
1500 997
1499 997
1499 1026
1 7 65 0 0 8320 0 84 94 0 0 3
1401 998
1403 998
1403 1025
1 7 66 0 0 8320 0 85 93 0 0 3
1306 993
1307 993
1307 1025
0 2 67 0 0 8320 0 0 87 103 0 5
1731 1248
1731 1262
1367 1262
1367 1228
1359 1228
0 1 2 0 0 0 0 0 87 78 0 3
1288 1205
1288 1228
1323 1228
1 0 68 0 0 4096 0 90 0 0 100 2
1787 1097
1787 1146
2 0 69 0 0 4096 0 90 0 0 101 2
1796 1097
1796 1134
3 0 70 0 0 4096 0 90 0 0 102 4
1805 1097
1805 1118
1806 1118
1806 1123
4 0 2 0 0 0 0 88 0 0 78 2
1718 1242
1718 1271
4 0 2 0 0 0 0 93 0 0 78 2
1352 1095
1352 1205
4 0 2 0 0 0 0 94 0 0 78 2
1448 1095
1448 1205
4 0 2 0 0 0 0 96 0 0 78 2
1544 1096
1544 1205
4 0 2 0 0 0 0 95 0 0 78 2
1640 1096
1640 1205
4 0 2 0 0 4096 0 90 0 0 78 2
1832 1097
1832 1271
4 0 2 0 0 0 0 92 0 0 78 2
1928 1097
1928 1271
1 4 2 0 0 4224 0 1 91 0 0 5
1255 1205
1644 1205
1644 1271
2023 1271
2023 1097
1 0 68 0 0 4096 0 93 0 0 100 2
1307 1095
1307 1146
2 0 69 0 0 4096 0 93 0 0 101 2
1316 1095
1316 1134
3 0 70 0 0 4096 0 93 0 0 102 2
1325 1095
1325 1123
1 0 68 0 0 0 0 94 0 0 100 4
1403 1095
1403 1141
1404 1141
1404 1146
2 0 69 0 0 0 0 94 0 0 101 2
1412 1095
1412 1134
3 0 70 0 0 0 0 94 0 0 102 2
1421 1095
1421 1123
1 0 68 0 0 0 0 96 0 0 100 2
1499 1096
1499 1146
2 0 69 0 0 0 0 96 0 0 101 2
1508 1096
1508 1134
3 0 70 0 0 0 0 96 0 0 102 2
1517 1096
1517 1123
1 0 68 0 0 0 0 95 0 0 100 2
1595 1096
1595 1146
2 0 69 0 0 0 0 95 0 0 101 2
1604 1096
1604 1134
3 0 70 0 0 0 0 95 0 0 102 2
1613 1096
1613 1123
1 0 68 0 0 0 0 89 0 0 100 2
1691 1096
1691 1146
2 0 69 0 0 0 0 89 0 0 101 2
1700 1096
1700 1134
3 0 70 0 0 0 0 89 0 0 102 2
1709 1096
1709 1123
1 0 68 0 0 0 0 92 0 0 100 2
1883 1097
1883 1146
2 0 69 0 0 0 0 92 0 0 101 2
1892 1097
1892 1134
3 0 70 0 0 0 0 92 0 0 102 2
1901 1097
1901 1123
1 1 71 0 0 8320 0 2 88 0 0 4
1120 1062
1120 1256
1673 1256
1673 1242
1 2 72 0 0 8320 0 7 88 0 0 4
1146 1064
1146 1251
1682 1251
1682 1242
1 3 73 0 0 8320 0 6 88 0 0 4
1178 1063
1178 1246
1691 1246
1691 1242
1 1 68 0 0 8320 0 3 91 0 0 4
1209 1062
1209 1146
1978 1146
1978 1097
1 2 69 0 0 8320 0 4 91 0 0 4
1233 1061
1233 1134
1987 1134
1987 1097
1 3 70 0 0 8320 0 5 91 0 0 4
1259 1060
1259 1123
1996 1123
1996 1097
5 6 67 0 0 0 0 88 88 0 0 2
1727 1248
1736 1248
5 0 74 0 0 8192 0 91 0 0 119 3
2032 1103
2032 1106
2041 1106
5 0 75 0 0 8192 0 92 0 0 118 3
1937 1103
1937 1106
1946 1106
5 0 76 0 0 8192 0 90 0 0 117 3
1841 1103
1841 1107
1850 1107
5 0 77 0 0 8192 0 89 0 0 116 3
1745 1102
1745 1105
1754 1105
6 0 78 0 0 8192 0 95 0 0 112 3
1658 1102
1658 1103
1649 1103
6 0 79 0 0 8192 0 96 0 0 113 3
1562 1102
1562 1104
1553 1104
6 0 80 0 0 8192 0 94 0 0 114 3
1466 1101
1466 1103
1457 1103
6 0 81 0 0 8192 0 93 0 0 115 3
1370 1101
1370 1104
1361 1104
10 5 78 0 0 12416 0 88 95 0 0 4
1700 1172
1700 1155
1649 1155
1649 1102
5 9 79 0 0 8320 0 96 88 0 0 4
1553 1102
1553 1160
1691 1160
1691 1172
5 8 80 0 0 8320 0 94 88 0 0 4
1457 1101
1457 1165
1682 1165
1682 1172
5 7 81 0 0 8320 0 93 88 0 0 3
1361 1101
1361 1172
1673 1172
6 11 77 0 0 4224 0 89 88 0 0 4
1754 1102
1754 1154
1709 1154
1709 1172
6 12 76 0 0 8320 0 90 88 0 0 4
1850 1103
1850 1159
1718 1159
1718 1172
6 13 75 0 0 8320 0 92 88 0 0 4
1946 1103
1946 1166
1727 1166
1727 1172
14 6 74 0 0 8320 0 88 91 0 0 4
1736 1172
1736 1171
2041 1171
2041 1103
1 14 82 0 0 8320 0 128 131 0 0 4
1897 441
1897 490
1663 490
1663 543
1 13 83 0 0 8320 0 127 131 0 0 4
1872 442
1872 500
1654 500
1654 543
1 12 84 0 0 8320 0 126 131 0 0 4
1845 441
1845 495
1645 495
1645 543
1 11 85 0 0 8320 0 125 131 0 0 4
1820 441
1820 515
1636 515
1636 543
1 10 86 0 0 8320 0 124 131 0 0 4
1796 443
1796 520
1627 520
1627 543
1 9 87 0 0 8320 0 123 131 0 0 4
1772 442
1772 525
1618 525
1618 543
1 8 88 0 0 8320 0 122 131 0 0 4
1746 443
1746 530
1609 530
1609 543
1 7 89 0 0 8320 0 121 131 0 0 4
1723 443
1723 535
1600 535
1600 543
1 14 90 0 0 8320 0 120 130 0 0 4
1697 444
1697 511
1563 511
1563 544
1 13 91 0 0 8320 0 119 130 0 0 4
1672 445
1672 505
1554 505
1554 544
1 12 92 0 0 8320 0 118 130 0 0 4
1646 446
1646 488
1545 488
1545 544
1 11 93 0 0 8320 0 117 130 0 0 4
1620 446
1620 484
1536 484
1536 544
1 10 94 0 0 8320 0 116 130 0 0 4
1596 446
1596 479
1527 479
1527 544
1 9 95 0 0 12416 0 115 130 0 0 4
1571 447
1571 475
1518 475
1518 544
1 8 96 0 0 12416 0 114 130 0 0 4
1546 447
1546 471
1509 471
1509 544
1 7 97 0 0 12416 0 113 130 0 0 4
1523 448
1523 467
1500 467
1500 544
1 14 98 0 0 12416 0 97 132 0 0 4
1504 448
1504 462
1429 462
1429 546
1 13 99 0 0 12416 0 98 132 0 0 4
1479 449
1479 458
1420 458
1420 546
1 12 100 0 0 12416 0 99 132 0 0 4
1452 448
1452 454
1411 454
1411 546
1 11 101 0 0 12416 0 100 132 0 0 4
1427 448
1427 452
1402 452
1402 546
1 10 102 0 0 8320 0 101 132 0 0 3
1403 450
1393 450
1393 546
1 9 103 0 0 4224 0 102 132 0 0 4
1379 449
1379 538
1384 538
1384 546
1 8 104 0 0 4224 0 103 132 0 0 4
1353 450
1353 503
1375 503
1375 546
1 7 105 0 0 4224 0 104 132 0 0 4
1330 450
1330 508
1366 508
1366 546
1 14 106 0 0 4224 0 105 133 0 0 4
1304 451
1304 503
1314 503
1314 546
1 13 107 0 0 4224 0 106 133 0 0 4
1279 452
1279 508
1305 508
1305 546
1 12 108 0 0 4224 0 107 133 0 0 4
1253 453
1253 513
1296 513
1296 546
1 11 109 0 0 4224 0 108 133 0 0 4
1227 453
1227 518
1287 518
1287 546
1 10 110 0 0 8320 0 109 133 0 0 4
1203 453
1203 523
1278 523
1278 546
1 9 111 0 0 8320 0 110 133 0 0 4
1178 454
1178 528
1269 528
1269 546
1 8 112 0 0 8320 0 111 133 0 0 4
1153 454
1153 533
1260 533
1260 546
1 7 113 0 0 8320 0 112 133 0 0 4
1130 455
1130 538
1251 538
1251 546
0 11 114 0 0 8320 0 0 129 169 0 4
1310 627
1310 664
1473 664
1473 682
0 12 115 0 0 8320 0 0 129 167 0 4
1424 626
1424 674
1482 674
1482 682
0 13 116 0 0 8320 0 0 129 168 0 4
1559 625
1559 664
1491 664
1491 682
0 14 117 0 0 8320 0 0 129 165 0 4
1659 624
1659 674
1500 674
1500 682
6 0 118 0 0 4096 0 129 0 0 158 2
1500 758
1500 757
5 0 118 0 0 0 0 129 0 0 158 2
1491 758
1491 757
1 1 118 0 0 8320 0 8 129 0 0 4
1784 651
1784 757
1437 757
1437 752
4 0 119 0 0 8192 0 129 0 0 166 4
1482 752
1482 772
1749 772
1749 669
1 2 120 0 0 8320 0 10 129 0 0 4
1030 608
1030 773
1446 773
1446 752
1 3 121 0 0 8320 0 11 129 0 0 4
1062 607
1062 763
1455 763
1455 752
4 0 119 0 0 0 0 132 0 0 166 2
1411 616
1411 669
4 0 119 0 0 0 0 130 0 0 166 2
1545 614
1545 669
4 0 119 0 0 0 0 131 0 0 166 2
1645 613
1645 669
5 6 117 0 0 0 0 131 131 0 0 4
1654 619
1654 624
1663 624
1663 619
4 1 119 0 0 8320 0 133 9 0 0 4
1296 616
1296 669
1749 669
1749 651
5 6 115 0 0 0 0 132 132 0 0 4
1420 622
1420 626
1429 626
1429 622
5 6 116 0 0 0 0 130 130 0 0 4
1554 620
1554 625
1563 625
1563 620
5 6 114 0 0 0 0 133 133 0 0 4
1305 622
1305 627
1314 627
1314 622
1 0 122 0 0 4096 0 130 0 0 176 2
1500 614
1500 660
1 0 122 0 0 0 0 132 0 0 176 2
1366 616
1366 660
1 0 122 0 0 0 0 133 0 0 176 2
1251 616
1251 660
2 0 123 0 0 4096 0 133 0 0 177 2
1260 616
1260 649
2 0 123 0 0 0 0 132 0 0 177 2
1375 616
1375 649
2 0 123 0 0 4096 0 130 0 0 177 2
1509 614
1509 649
1 1 122 0 0 8320 0 14 131 0 0 4
1093 606
1093 660
1600 660
1600 613
1 2 123 0 0 8320 0 13 131 0 0 4
1117 605
1117 649
1609 649
1609 613
3 0 124 0 0 4096 0 133 0 0 181 2
1269 616
1269 638
3 0 124 0 0 0 0 132 0 0 181 2
1384 616
1384 638
3 0 124 0 0 4096 0 130 0 0 181 2
1518 614
1518 638
1 3 124 0 0 8320 0 12 131 0 0 4
1143 604
1143 638
1618 638
1618 613
1 1 125 0 0 8320 0 17 142 0 0 3
120 590
120 665
442 665
1 2 126 0 0 8320 0 18 142 0 0 3
150 591
150 674
442 674
1 3 127 0 0 8320 0 19 142 0 0 3
179 594
179 683
442 683
0 6 128 0 0 4096 0 0 142 186 0 2
395 728
436 728
1 5 128 0 0 4224 0 15 142 0 0 4
131 794
395 794
395 719
436 719
1 4 129 0 0 4224 0 16 142 0 0 4
131 766
323 766
323 710
442 710
7 1 130 0 0 4224 0 142 141 0 0 3
512 665
588 665
588 631
8 1 131 0 0 4224 0 142 140 0 0 3
512 674
611 674
611 630
9 1 132 0 0 4224 0 142 139 0 0 3
512 683
636 683
636 630
10 1 133 0 0 4224 0 142 138 0 0 3
512 692
661 692
661 629
11 1 134 0 0 4224 0 142 137 0 0 3
512 701
685 701
685 629
12 1 135 0 0 4224 0 142 136 0 0 3
512 710
707 710
707 627
13 1 136 0 0 4224 0 142 135 0 0 3
512 719
736 719
736 625
14 1 137 0 0 4224 0 142 134 0 0 3
512 728
762 728
762 625
2 0 138 0 0 8192 0 143 0 0 197 4
191 223
281 223
281 334
286 334
1 1 138 0 0 4224 0 144 152 0 0 4
446 345
286 345
286 318
445 318
0 0 139 0 0 4096 0 0 0 200 199 4
109 196
303 196
303 213
308 213
1 1 139 0 0 0 0 145 153 0 0 4
453 237
308 237
308 212
453 212
0 1 139 0 0 0 0 0 143 207 0 3
109 61
109 223
155 223
1 0 140 0 0 8192 0 21 0 0 202 4
90 116
102 116
102 306
230 306
3 3 140 0 0 12416 0 157 156 0 0 4
591 260
230 260
230 363
595 363
0 0 140 0 0 0 0 0 0 206 204 4
142 95
322 95
322 136
449 136
1 1 140 0 0 0 0 146 154 0 0 4
457 150
449 150
449 120
457 120
3 0 139 0 0 4224 0 158 0 0 207 3
590 171
190 171
190 53
1 1 140 0 0 0 0 21 155 0 0 4
90 116
142 116
142 27
458 27
1 1 139 0 0 0 0 22 147 0 0 4
91 61
164 61
164 53
457 53
1 3 141 0 0 4224 0 20 159 0 0 4
487 80
576 80
576 79
584 79
4 1 142 0 0 4224 0 156 148 0 0 3
640 354
780 354
780 342
4 1 143 0 0 12416 0 157 149 0 0 5
636 251
709 251
709 252
784 252
784 249
4 1 144 0 0 4224 0 158 150 0 0 3
635 162
779 162
779 156
4 1 145 0 0 4224 0 159 151 0 0 3
629 70
779 70
779 65
2 2 146 0 0 4224 0 144 156 0 0 4
482 345
587 345
587 354
595 354
2 2 147 0 0 4224 0 145 157 0 0 4
489 237
583 237
583 251
591 251
2 2 148 0 0 12416 0 146 158 0 0 4
493 150
541 150
541 162
590 162
2 2 149 0 0 4224 0 147 159 0 0 4
493 53
540 53
540 70
584 70
2 1 150 0 0 4224 0 152 156 0 0 4
481 318
580 318
580 345
595 345
2 1 151 0 0 4224 0 153 157 0 0 4
489 212
576 212
576 242
591 242
1 2 152 0 0 12416 0 158 154 0 0 4
590 153
555 153
555 120
493 120
2 1 153 0 0 12416 0 155 159 0 0 4
494 27
519 27
519 61
584 61
96
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1110 385 1145 406
1119 392 1135 407
2 31
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1140 384 1173 405
1148 391 1164 406
2 30
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1163 384 1198 405
1172 391 1188 406
2 29
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1189 382 1224 403
1198 389 1214 404
2 28
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1213 387 1248 408
1222 393 1238 408
2 27
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1237 384 1270 405
1245 391 1261 406
2 26
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1262 383 1295 404
1270 390 1286 405
2 25
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1291 383 1324 404
1299 389 1315 404
2 24
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1317 383 1352 404
1326 389 1342 404
2 23
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1339 385 1372 406
1347 392 1363 407
2 22
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1362 380 1397 401
1371 387 1387 402
2 21
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1386 385 1419 406
1394 392 1410 407
2 20
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1414 383 1447 404
1422 390 1438 405
2 19
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1437 385 1472 406
1446 392 1462 407
2 18
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1463 381 1498 402
1472 388 1488 403
2 17
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1487 381 1522 402
1496 388 1512 403
2 16
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1507 381 1542 402
1516 387 1532 402
2 15
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1529 381 1562 402
1537 388 1553 403
2 14
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1555 379 1590 400
1564 386 1580 401
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1579 380 1614 401
1588 387 1604 402
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1604 381 1639 402
1613 387 1629 402
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1630 380 1663 401
1638 386 1654 401
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1661 376 1686 397
1669 383 1677 398
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1684 376 1711 397
1693 383 1701 398
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1710 382 1737 403
1719 388 1727 403
1 7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1733 380 1760 401
1742 386 1750 401
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1759 377 1786 398
1768 384 1776 399
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1780 378 1805 399
1788 385 1796 400
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1807 376 1834 397
1816 383 1824 398
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1828 376 1855 397
1837 383 1845 398
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1857 376 1884 397
1866 382 1874 397
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1884 379 1911 400
1893 385 1901 400
1 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1973 807 2000 828
1982 813 1990 828
1 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1973 833 2000 854
1982 839 1990 854
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1976 857 2003 878
1985 864 1993 879
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1975 875 2002 896
1984 882 1992 897
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1973 898 1998 919
1981 905 1989 920
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1970 924 1997 945
1979 931 1987 946
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1970 943 1997 964
1979 949 1987 964
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1967 965 1994 986
1976 971 1984 986
1 7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1876 823 1903 844
1885 830 1893 845
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1881 845 1906 866
1889 852 1897 867
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1876 865 1911 886
1885 872 1901 887
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1875 887 1908 908
1883 894 1899 909
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1876 907 1909 928
1884 913 1900 928
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1876 931 1911 952
1885 938 1901 953
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1872 955 1905 976
1880 961 1896 976
2 14
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1871 975 1904 996
1879 981 1895 996
2 15
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1769 820 1804 841
1778 827 1794 842
2 16
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1770 846 1803 867
1778 852 1794 867
2 17
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1772 865 1805 886
1780 872 1796 887
2 18
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1775 888 1808 909
1783 895 1799 910
2 19
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1771 908 1806 929
1780 915 1796 930
2 20
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1775 930 1810 951
1784 937 1800 952
2 21
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1774 954 1809 975
1783 961 1799 976
2 22
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1773 975 1806 996
1781 982 1797 997
2 23
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1676 810 1709 831
1684 817 1700 832
2 24
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1678 837 1711 858
1686 844 1702 859
2 25
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1680 859 1713 880
1688 866 1704 881
2 26
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1679 880 1714 901
1688 886 1704 901
2 27
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1677 904 1712 925
1686 911 1702 926
2 28
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1676 926 1711 947
1685 933 1701 948
2 29
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1678 946 1711 967
1686 953 1702 968
2 30
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1673 972 1708 993
1682 979 1698 994
2 31
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1585 819 1620 840
1594 825 1610 840
2 32
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1584 840 1617 861
1592 847 1608 862
2 33
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1583 863 1618 884
1592 869 1608 884
2 34
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1583 881 1616 902
1591 888 1607 903
2 35
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1583 905 1616 926
1591 912 1607 927
2 36
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1584 927 1617 948
1592 934 1608 949
2 37
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1583 947 1616 968
1591 954 1607 969
2 38
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1579 971 1612 992
1587 978 1603 993
2 39
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1490 819 1523 840
1498 825 1514 840
2 40
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1486 840 1521 861
1495 847 1511 862
2 41
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1488 863 1523 884
1497 870 1513 885
2 42
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1490 884 1523 905
1498 890 1514 905
2 43
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1488 909 1521 930
1496 916 1512 931
2 44
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1488 930 1521 951
1496 937 1512 952
2 45
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1485 951 1518 972
1493 958 1509 973
2 46
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1484 975 1517 996
1492 982 1508 997
2 47
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1391 815 1426 836
1400 822 1416 837
2 48
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1391 839 1424 860
1399 846 1415 861
2 49
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1397 858 1430 879
1405 864 1421 879
2 50
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1397 876 1432 897
1406 883 1422 898
2 51
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1395 904 1428 925
1403 911 1419 926
2 52
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1395 925 1428 946
1403 931 1419 946
2 53
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1389 948 1424 969
1398 954 1414 969
2 54
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1386 974 1421 995
1395 981 1411 996
2 55
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1297 815 1330 836
1305 822 1321 837
2 56
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1294 841 1329 862
1303 847 1319 862
2 57
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1298 859 1331 880
1306 866 1322 881
2 58
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1299 879 1332 900
1307 885 1323 900
2 59
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1294 904 1329 925
1303 910 1319 925
2 60
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1293 926 1328 947
1302 933 1318 948
2 61
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1294 944 1327 965
1302 951 1318 966
2 62
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1289 973 1324 994
1298 980 1314 995
2 63
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
