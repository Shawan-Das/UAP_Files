CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 930 1 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
61
13 Logic Switch~
5 370 1285 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3805 0 0
2
44291.8 0
0
13 Logic Switch~
5 287 929 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
7 Control
-68 -4 -19 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5219 0 0
2
44291.8 1
0
13 Logic Switch~
5 317 840 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3795 0 0
2
44291.8 2
0
13 Logic Switch~
5 602 441 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3637 0 0
2
44291.8 3
0
13 Logic Switch~
5 135 473 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3226 0 0
2
44291.8 4
0
13 Logic Switch~
5 556 142 0 1 11
0 37
0
0 0 21360 90
2 0V
-8 13 6 21
7 Control
-38 26 11 34
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6966 0 0
2
44291.8 5
0
13 Logic Switch~
5 579 214 0 1 11
0 44
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9796 0 0
2
44291.8 6
0
13 Logic Switch~
5 359 225 0 1 11
0 52
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5952 0 0
2
44291.8 7
0
13 Logic Switch~
5 156 226 0 1 11
0 54
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3649 0 0
2
44291.8 8
0
12 Hex Display~
7 553 767 0 18 19
10 15 14 13 59 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP4
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
3716 0 0
2
5.8998e-315 0
0
12 Hex Display~
7 884 368 0 18 19
10 21 22 23 60 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
4797 0 0
2
5.8998e-315 0
0
12 Hex Display~
7 765 1064 0 16 19
10 4 3 2 61 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
4681 0 0
2
5.8998e-315 0
0
8 2-In OR~
219 552 1272 0 3 22
0 4 6 8
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U15A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
9730 0 0
2
5.8998e-315 0
0
9 2-In AND~
219 492 1135 0 3 22
0 3 2 10
0
0 0 624 180
5 74F08
-18 -24 17 -16
4 U14A
-15 -4 13 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
9874 0 0
2
5.8998e-315 0
0
9 2-In AND~
219 733 1163 0 3 22
0 5 3 7
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7D
-11 0 10 8
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
364 0 0
2
5.8998e-315 0
0
5 4027~
219 489 1238 0 7 32
0 62 10 9 11 63 5 4
0
0 0 4720 0
4 4027
7 -60 35 -52
4 U13B
6 -63 34 -55
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 10 0
1 U
3656 0 0
2
44291.8 9
0
5 4027~
219 642 1238 0 7 32
0 64 5 9 8 65 66 3
0
0 0 4720 0
4 4027
7 -60 35 -52
4 U13A
-31 -60 -3 -52
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 10 0
1 U
3131 0 0
2
44291.8 10
0
5 4027~
219 812 1238 0 7 32
0 67 7 9 4 68 6 2
0
0 0 4720 0
4 4027
7 -60 35 -52
4 U10B
4 -62 32 -54
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 8 0
1 U
6772 0 0
2
44291.8 11
0
7 Pulser~
4 328 1208 0 10 12
0 9 69 9 70 0 0 5 5 3
8
0
0 0 4656 270
0
3 V17
-40 -3 -19 5
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9557 0 0
2
44291.8 12
0
14 Logic Display~
6 644 1079 0 1 2
10 71
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L21
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
5789 0 0
2
44291.8 13
0
14 Logic Display~
6 665 1079 0 1 2
10 72
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L20
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
7328 0 0
2
44291.8 14
0
14 Logic Display~
6 686 1080 0 1 2
10 73
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
4799 0 0
2
44291.8 15
0
9 2-In XOR~
219 494 861 0 3 22
0 15 12 16
0
0 0 624 0
5 74F86
-18 -24 17 -16
4 U12A
-494 -836 -466 -828
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
9196 0 0
2
44291.8 16
0
9 2-In XOR~
219 682 860 0 3 22
0 14 12 18
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U4D
40 -347 61 -339
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3857 0 0
2
44291.8 17
0
9 2-In AND~
219 745 832 0 3 22
0 16 18 17
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7C
-15 -5 6 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
7125 0 0
2
44291.8 18
0
7 Pulser~
4 259 858 0 10 12
0 20 74 20 75 0 0 5 5 3
8
0
0 0 4656 270
0
3 V15
-40 -3 -19 5
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3641 0 0
2
44291.8 19
0
5 4027~
219 802 884 0 7 32
0 76 17 20 17 77 78 13
0
0 0 4720 0
4 4027
7 -60 35 -52
4 U10A
4 -62 32 -54
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 8 0
1 U
9821 0 0
2
44291.8 20
0
5 4027~
219 620 887 0 7 32
0 79 16 20 16 80 81 14
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U9B
-28 -60 -7 -52
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 7 0
1 U
3187 0 0
2
44291.8 21
0
5 4027~
219 420 888 0 7 32
0 82 19 20 19 83 84 15
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U9A
3 -60 24 -52
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 7 0
1 U
762 0 0
2
44291.8 22
0
5 4027~
219 710 518 0 7 32
0 29 27 30 27 85 26 21
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U8B
3 -60 24 -52
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 6 0
1 U
39 0 0
2
44291.8 23
0
5 4027~
219 798 516 0 7 32
0 86 26 30 26 28 25 22
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U8A
-28 -60 -7 -52
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 6 0
1 U
9450 0 0
2
44291.8 24
0
5 4027~
219 887 515 0 7 32
0 87 24 30 24 88 89 23
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U6B
7 -62 28 -54
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 4 0
1 U
3236 0 0
2
44291.8 25
0
7 Pulser~
4 549 488 0 10 12
0 30 90 30 91 0 0 5 5 3
8
0
0 0 4656 270
0
3 V12
-40 -3 -19 5
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3321 0 0
2
44291.8 26
0
9 2-In AND~
219 849 427 0 3 22
0 26 25 24
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7B
-12 -2 9 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
8879 0 0
2
44291.8 27
0
9 2-In AND~
219 383 456 0 3 22
0 31 32 34
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
5433 0 0
2
44291.8 28
0
7 Pulser~
4 82 520 0 10 12
0 36 92 36 93 0 0 5 5 3
8
0
0 0 4656 270
0
2 V8
-37 -3 -23 5
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3679 0 0
2
44291.8 29
0
5 4027~
219 420 547 0 7 32
0 94 34 36 34 95 96 33
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U6A
7 -62 28 -54
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 4 0
1 U
9342 0 0
2
44291.8 30
0
5 4027~
219 331 548 0 7 32
0 97 31 36 31 98 99 32
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U5B
-28 -60 -7 -52
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 3 0
1 U
3623 0 0
2
44291.8 31
0
5 4027~
219 243 550 0 7 32
0 100 35 36 35 101 102 31
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U5A
3 -60 24 -52
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 3 0
1 U
3722 0 0
2
44291.8 32
0
9 2-In XOR~
219 701 95 0 3 22
0 37 39 40
0
0 0 624 90
5 74F86
-18 -24 17 -16
3 U4C
-81 -385 -60 -377
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
8993 0 0
2
44291.8 33
0
9 2-In XOR~
219 655 93 0 3 22
0 37 43 42
0
0 0 624 90
5 74F86
-18 -24 17 -16
3 U4B
-83 -351 -62 -343
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3723 0 0
2
44291.8 34
0
9 2-In XOR~
219 600 95 0 3 22
0 37 38 41
0
0 0 624 90
5 74F86
-18 -24 17 -16
3 U4A
-79 -310 -58 -302
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
6244 0 0
2
44291.8 35
0
7 74LS293
154 668 167 0 8 17
0 44 44 103 45 38 43 39 104
0
0 0 4848 90
7 74LS293
-24 -35 25 -27
2 U3
30 -7 44 1
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 512 1 0 0 0
1 U
6421 0 0
2
44291.8 36
0
7 Pulser~
4 662 261 0 10 12
0 45 105 45 106 0 0 5 5 3
8
0
0 0 4656 0
0
2 V6
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7743 0 0
2
44291.8 37
0
14 Logic Display~
6 688 35 0 1 2
10 40
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9840 0 0
2
44291.8 38
0
14 Logic Display~
6 658 35 0 1 2
10 42
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6910 0 0
2
44291.8 39
0
14 Logic Display~
6 626 35 0 1 2
10 41
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
449 0 0
2
44291.8 40
0
9 Inverter~
13 463 110 0 2 22
0 47 49
0
0 0 624 90
5 74F04
-18 -19 17 -11
3 U2C
-463 -88 -442 -80
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
8761 0 0
2
44291.8 41
0
9 Inverter~
13 441 110 0 2 22
0 48 50
0
0 0 624 90
5 74F04
-18 -19 17 -11
3 U2B
-439 -106 -418 -98
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
6748 0 0
2
44291.8 42
0
9 Inverter~
13 420 110 0 2 22
0 46 51
0
0 0 624 90
5 74F04
-18 -19 17 -11
3 U2A
-420 -96 -399 -88
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
7393 0 0
2
44291.8 43
0
7 74LS293
154 448 178 0 8 17
0 52 52 107 53 46 48 47 108
0
0 0 4848 90
7 74LS293
-24 -35 25 -27
2 U1
30 -7 44 1
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 512 1 0 0 0
1 U
7699 0 0
2
44291.8 44
0
7 Pulser~
4 442 272 0 10 12
0 53 109 53 110 0 0 5 5 3
8
0
0 0 4656 0
0
2 V4
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6638 0 0
2
44291.8 45
0
14 Logic Display~
6 465 62 0 1 2
10 49
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4595 0 0
2
44291.8 46
0
14 Logic Display~
6 444 61 0 1 2
10 50
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9395 0 0
2
44291.8 47
0
14 Logic Display~
6 423 61 0 1 2
10 51
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3303 0 0
2
44291.8 48
0
14 Logic Display~
6 220 62 0 1 2
10 55
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4498 0 0
2
44291.8 49
0
14 Logic Display~
6 241 62 0 1 2
10 56
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9728 0 0
2
44291.8 50
0
14 Logic Display~
6 262 61 0 1 2
10 57
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3789 0 0
2
44291.8 51
0
12 Hex Display~
7 418 384 0 18 19
10 31 32 33 111 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
3978 0 0
2
44291.8 52
0
7 Pulser~
4 239 273 0 10 12
0 58 112 58 113 0 0 5 5 3
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3494 0 0
2
44291.8 53
0
7 74LS293
154 245 179 0 8 17
0 54 54 114 58 55 56 57 115
0
0 0 4848 90
7 74LS293
-24 -35 25 -27
3 U11
27 -7 48 1
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 512 1 0 0 0
1 U
3507 0 0
2
44291.8 54
0
100
3 0 2 0 0 4096 0 12 0 0 4 2
762 1088
762 1126
0 2 3 0 0 4096 0 0 12 5 0 3
676 1146
768 1146
768 1088
0 1 4 0 0 4112 0 0 12 7 0 4
758 1249
758 1213
774 1213
774 1088
7 2 2 0 0 12416 0 18 14 0 0 4
836 1202
846 1202
846 1126
510 1126
0 1 3 0 0 12416 0 0 14 9 0 4
701 1180
676 1180
676 1144
510 1144
2 0 5 0 0 4096 0 17 0 0 8 4
618 1202
609 1202
609 1203
604 1203
0 4 4 0 0 4224 0 0 18 11 0 4
531 1249
775 1249
775 1220
788 1220
6 1 5 0 0 12416 0 16 15 0 0 4
519 1220
604 1220
604 1154
709 1154
7 2 3 0 0 0 0 17 15 0 0 4
666 1202
701 1202
701 1172
709 1172
6 2 6 0 0 12416 0 18 13 0 0 6
842 1220
846 1220
846 1292
531 1292
531 1281
539 1281
7 1 4 0 0 0 0 16 13 0 0 4
513 1202
531 1202
531 1263
539 1263
3 2 7 0 0 8320 0 15 18 0 0 4
754 1163
780 1163
780 1202
788 1202
3 4 8 0 0 8320 0 13 17 0 0 4
585 1272
610 1272
610 1220
618 1220
3 0 9 0 0 8192 0 17 0 0 15 3
618 1211
614 1211
614 1302
0 3 9 0 0 12416 0 0 18 18 0 6
428 1211
427 1211
427 1302
780 1302
780 1211
788 1211
3 2 10 0 0 8320 0 14 16 0 0 4
465 1135
457 1135
457 1202
465 1202
1 4 11 0 0 12416 0 1 16 0 0 4
382 1285
394 1285
394 1220
465 1220
0 3 9 0 0 0 0 0 16 19 0 2
351 1211
465 1211
1 3 9 0 0 0 0 19 19 0 0 6
336 1185
336 1184
351 1184
351 1235
336 1235
336 1233
1 0 12 0 0 4096 0 2 0 0 24 2
299 929
457 929
7 3 13 0 0 12416 0 27 10 0 0 5
826 848
836 848
836 812
550 812
550 791
0 2 14 0 0 8320 0 0 10 29 0 4
654 851
654 807
556 807
556 791
0 1 15 0 0 8320 0 0 10 30 0 4
458 852
458 834
562 834
562 791
2 2 12 0 0 12416 0 23 24 0 0 6
478 870
457 870
457 929
658 929
658 869
666 869
0 1 16 0 0 8320 0 0 25 26 0 3
569 844
569 823
721 823
3 0 16 0 0 0 0 23 0 0 32 5
527 861
532 861
532 844
569 844
569 851
3 0 17 0 0 8320 0 25 0 0 31 4
766 832
771 832
771 851
770 851
2 3 18 0 0 8320 0 25 24 0 0 4
721 841
714 841
714 860
715 860
7 1 14 0 0 0 0 28 24 0 0 2
644 851
666 851
7 1 15 0 0 0 0 29 23 0 0 2
444 852
478 852
2 4 17 0 0 0 0 27 27 0 0 4
778 848
770 848
770 866
778 866
2 4 16 0 0 0 0 28 28 0 0 4
596 851
569 851
569 869
596 869
1 0 19 0 0 4224 0 3 0 0 34 3
329 840
388 840
388 852
2 4 19 0 0 0 0 29 29 0 0 4
396 852
388 852
388 870
396 870
3 0 20 0 0 12416 0 27 0 0 37 5
778 857
761 857
761 907
312 907
312 861
3 0 20 0 0 0 0 28 0 0 35 3
596 860
561 860
561 907
0 3 20 0 0 0 0 0 29 38 0 2
282 861
396 861
1 3 20 0 0 0 0 26 26 0 0 6
267 835
267 834
282 834
282 885
267 885
267 883
7 1 21 0 0 12416 0 30 11 0 0 5
734 482
757 482
757 408
893 408
893 392
7 2 22 0 0 16512 0 31 11 0 0 5
822 480
843 480
843 449
887 449
887 392
7 3 23 0 0 8320 0 32 11 0 0 5
911 479
921 479
921 428
881 428
881 392
3 0 24 0 0 16512 0 34 0 0 46 5
870 427
873 427
873 444
855 444
855 479
6 2 25 0 0 8320 0 31 34 0 0 6
828 498
832 498
832 448
805 448
805 436
825 436
0 1 26 0 0 4224 0 0 34 45 0 3
747 500
747 418
825 418
6 0 26 0 0 0 0 30 0 0 47 4
740 500
761 500
761 498
766 498
2 4 24 0 0 0 0 32 32 0 0 4
863 479
855 479
855 497
863 497
2 4 26 0 0 0 0 31 31 0 0 4
774 480
766 480
766 498
774 498
1 0 27 0 0 4224 0 4 0 0 49 3
614 441
678 441
678 482
2 4 27 0 0 0 0 30 30 0 0 4
686 482
678 482
678 500
686 500
5 0 28 0 0 4224 0 31 0 0 0 2
798 522
798 527
1 0 29 0 0 4224 0 30 0 0 0 2
710 461
710 455
3 0 30 0 0 12416 0 32 0 0 54 5
863 488
846 488
846 544
602 544
602 491
3 0 30 0 0 0 0 31 0 0 52 3
774 489
755 489
755 544
0 3 30 0 0 0 0 0 30 55 0 2
572 491
686 491
1 3 30 0 0 0 0 33 33 0 0 6
557 465
557 464
572 464
572 515
557 515
557 513
0 1 31 0 0 8320 0 0 59 59 0 4
338 437
338 427
427 427
427 408
0 2 32 0 0 12416 0 0 59 60 0 4
369 481
369 480
421 480
421 408
7 3 33 0 0 8320 0 37 59 0 0 5
444 511
454 511
454 445
415 445
415 408
0 1 31 0 0 0 0 0 35 62 0 5
280 514
280 437
338 437
338 447
359 447
7 2 32 0 0 0 0 38 35 0 0 6
355 512
369 512
369 481
352 481
352 465
359 465
3 0 34 0 0 16512 0 35 0 0 63 5
404 456
408 456
408 476
391 476
391 511
7 0 31 0 0 0 0 39 0 0 64 3
267 514
299 514
299 512
2 4 34 0 0 0 0 37 37 0 0 4
396 511
388 511
388 529
396 529
2 4 31 0 0 0 0 38 38 0 0 4
307 512
299 512
299 530
307 530
1 0 35 0 0 4224 0 5 0 0 66 3
147 473
211 473
211 514
2 4 35 0 0 0 0 39 39 0 0 4
219 514
211 514
211 532
219 532
3 0 36 0 0 12416 0 37 0 0 69 5
396 520
379 520
379 576
135 576
135 523
3 0 36 0 0 0 0 38 0 0 67 3
307 521
288 521
288 576
0 3 36 0 0 0 0 0 39 70 0 2
105 523
219 523
1 3 36 0 0 0 0 36 36 0 0 6
90 497
90 496
105 496
105 547
90 547
90 545
1 0 37 0 0 4096 0 41 0 0 72 2
649 112
649 123
1 0 37 0 0 8320 0 40 0 0 73 3
695 114
695 123
594 123
1 1 37 0 0 0 0 6 42 0 0 4
557 129
557 128
594 128
594 114
5 2 38 0 0 8320 0 43 42 0 0 4
655 133
655 129
612 129
612 114
7 2 39 0 0 8320 0 43 40 0 0 4
673 133
673 129
713 129
713 114
3 1 40 0 0 8320 0 40 45 0 0 4
704 65
704 58
688 58
688 53
3 1 41 0 0 8320 0 42 47 0 0 4
603 65
603 60
626 60
626 53
3 1 42 0 0 4224 0 41 46 0 0 2
658 63
658 53
6 2 43 0 0 12416 0 43 41 0 0 4
664 133
664 125
667 125
667 112
1 0 44 0 0 4224 0 7 0 0 81 2
591 214
655 214
1 2 44 0 0 0 0 43 43 0 0 4
655 197
655 216
664 216
664 197
4 0 45 0 0 4096 0 43 0 0 83 2
682 203
682 238
1 3 45 0 0 12416 0 44 44 0 0 6
638 252
628 252
628 238
699 238
699 252
686 252
5 1 46 0 0 8320 0 51 50 0 0 4
435 144
435 136
423 136
423 128
7 1 47 0 0 8320 0 51 48 0 0 4
453 144
453 136
466 136
466 128
6 1 48 0 0 4224 0 51 49 0 0 2
444 144
444 128
1 2 49 0 0 12416 0 53 48 0 0 4
465 80
465 84
466 84
466 92
1 2 50 0 0 4224 0 54 49 0 0 2
444 79
444 92
1 2 51 0 0 4224 0 55 50 0 0 2
423 79
423 92
1 0 52 0 0 4224 0 8 0 0 91 2
371 225
435 225
1 2 52 0 0 0 0 51 51 0 0 4
435 208
435 227
444 227
444 208
4 0 53 0 0 4096 0 51 0 0 93 2
462 214
462 249
1 3 53 0 0 12416 0 52 52 0 0 6
418 263
408 263
408 249
480 249
480 263
466 263
1 0 54 0 0 4224 0 9 0 0 98 2
168 226
232 226
1 5 55 0 0 4224 0 56 61 0 0 4
220 80
220 118
232 118
232 145
1 6 56 0 0 4224 0 57 61 0 0 2
241 80
241 145
1 7 57 0 0 4224 0 58 61 0 0 4
262 79
262 117
250 117
250 145
1 2 54 0 0 0 0 61 61 0 0 4
232 209
232 228
241 228
241 209
4 0 58 0 0 4096 0 61 0 0 100 2
259 215
259 250
1 3 58 0 0 12416 0 60 60 0 0 6
215 264
205 264
205 250
277 250
277 264
263 264
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
162 294 309 315
171 300 299 315
16 MOD-8 Up-counter
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
363 294 524 315
371 300 515 315
18 Mod-8 Down-Counter
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
574 292 761 313
583 299 751 314
21 Mod-8 Up-Down Counter
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
207 579 354 600
216 585 344 600
16 MOD-8 Up-counter
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
691 549 852 570
699 555 843 570
18 Mod-8 Down-Counter
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
471 936 658 957
480 943 648 958
21 Mod-8 Up-Down Counter
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
